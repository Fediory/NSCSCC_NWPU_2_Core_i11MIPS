module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  reg  state_5; // @[PRNG.scala 55:49]
  reg  state_6; // @[PRNG.scala 55:49]
  reg  state_7; // @[PRNG.scala 55:49]
  reg  state_8; // @[PRNG.scala 55:49]
  reg  state_9; // @[PRNG.scala 55:49]
  reg  state_10; // @[PRNG.scala 55:49]
  reg  state_11; // @[PRNG.scala 55:49]
  reg  state_12; // @[PRNG.scala 55:49]
  reg  state_13; // @[PRNG.scala 55:49]
  reg  state_14; // @[PRNG.scala 55:49]
  reg  state_15; // @[PRNG.scala 55:49]
  wire  _T_2 = state_15 ^ state_13 ^ state_12 ^ state_10; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  assign io_out_5 = state_5; // @[PRNG.scala 78:10]
  assign io_out_6 = state_6; // @[PRNG.scala 78:10]
  assign io_out_7 = state_7; // @[PRNG.scala 78:10]
  assign io_out_8 = state_8; // @[PRNG.scala 78:10]
  assign io_out_9 = state_9; // @[PRNG.scala 78:10]
  assign io_out_10 = state_10; // @[PRNG.scala 78:10]
  assign io_out_11 = state_11; // @[PRNG.scala 78:10]
  assign io_out_12 = state_12; // @[PRNG.scala 78:10]
  assign io_out_13 = state_13; // @[PRNG.scala 78:10]
  assign io_out_14 = state_14; // @[PRNG.scala 78:10]
  assign io_out_15 = state_15; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T_2; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_4 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_4 <= state_3;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_5 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_5 <= state_4;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_6 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_6 <= state_5;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_7 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_7 <= state_6;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_8 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_8 <= state_7;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_9 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_9 <= state_8;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_10 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_10 <= state_9;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_11 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_11 <= state_10;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_12 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_12 <= state_11;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_13 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_13 <= state_12;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_14 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_14 <= state_13;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_15 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_15 <= state_14;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module dcache(
  input          clock,
  input          reset,
  input          valid,
  input          op,
  input  [7:0]   index,
  input  [19:0]  tag,
  input  [3:0]   offset,
  input  [3:0]   wstrb,
  input  [31:0]  wdata,
  output         addr_ok,
  output         data_ok,
  output [31:0]  rdata,
  input  [2:0]   lstype,
  input          uncached,
  output         rd_req,
  output [2:0]   rd_type,
  output [31:0]  rd_addr,
  input          rd_rdy,
  input          ret_valid,
  input          ret_last,
  input  [31:0]  ret_data,
  output         wr_req,
  output [2:0]   wr_type,
  output [31:0]  wr_addr,
  output [3:0]   wr_wstrb,
  output [127:0] wr_data,
  input          wr_rdy,
  input          cache_op_en,
  input  [2:0]   cache_op,
  input  [19:0]  cache_tag,
  input  [7:0]   cache_index,
  input  [3:0]   cache_offset,
  input  [21:0]  tag_input,
  output [21:0]  tag_output,
  output         cache_op_done,
  output         hit
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] tagv_ram_addra; // @[dcache.scala 110:49]
  wire  tagv_ram_clka; // @[dcache.scala 110:49]
  wire [20:0] tagv_ram_dina; // @[dcache.scala 110:49]
  wire [20:0] tagv_ram_douta; // @[dcache.scala 110:49]
  wire  tagv_ram_wea; // @[dcache.scala 110:49]
  wire [7:0] tagv_ram_1_addra; // @[dcache.scala 110:49]
  wire  tagv_ram_1_clka; // @[dcache.scala 110:49]
  wire [20:0] tagv_ram_1_dina; // @[dcache.scala 110:49]
  wire [20:0] tagv_ram_1_douta; // @[dcache.scala 110:49]
  wire  tagv_ram_1_wea; // @[dcache.scala 110:49]
  wire [7:0] data_ram_addra; // @[dcache.scala 111:65]
  wire  data_ram_clka; // @[dcache.scala 111:65]
  wire [31:0] data_ram_dina; // @[dcache.scala 111:65]
  wire [31:0] data_ram_douta; // @[dcache.scala 111:65]
  wire [3:0] data_ram_wea; // @[dcache.scala 111:65]
  wire [7:0] data_ram_1_addra; // @[dcache.scala 111:65]
  wire  data_ram_1_clka; // @[dcache.scala 111:65]
  wire [31:0] data_ram_1_dina; // @[dcache.scala 111:65]
  wire [31:0] data_ram_1_douta; // @[dcache.scala 111:65]
  wire [3:0] data_ram_1_wea; // @[dcache.scala 111:65]
  wire [7:0] data_ram_2_addra; // @[dcache.scala 111:65]
  wire  data_ram_2_clka; // @[dcache.scala 111:65]
  wire [31:0] data_ram_2_dina; // @[dcache.scala 111:65]
  wire [31:0] data_ram_2_douta; // @[dcache.scala 111:65]
  wire [3:0] data_ram_2_wea; // @[dcache.scala 111:65]
  wire [7:0] data_ram_3_addra; // @[dcache.scala 111:65]
  wire  data_ram_3_clka; // @[dcache.scala 111:65]
  wire [31:0] data_ram_3_dina; // @[dcache.scala 111:65]
  wire [31:0] data_ram_3_douta; // @[dcache.scala 111:65]
  wire [3:0] data_ram_3_wea; // @[dcache.scala 111:65]
  wire [7:0] data_ram_4_addra; // @[dcache.scala 111:65]
  wire  data_ram_4_clka; // @[dcache.scala 111:65]
  wire [31:0] data_ram_4_dina; // @[dcache.scala 111:65]
  wire [31:0] data_ram_4_douta; // @[dcache.scala 111:65]
  wire [3:0] data_ram_4_wea; // @[dcache.scala 111:65]
  wire [7:0] data_ram_5_addra; // @[dcache.scala 111:65]
  wire  data_ram_5_clka; // @[dcache.scala 111:65]
  wire [31:0] data_ram_5_dina; // @[dcache.scala 111:65]
  wire [31:0] data_ram_5_douta; // @[dcache.scala 111:65]
  wire [3:0] data_ram_5_wea; // @[dcache.scala 111:65]
  wire [7:0] data_ram_6_addra; // @[dcache.scala 111:65]
  wire  data_ram_6_clka; // @[dcache.scala 111:65]
  wire [31:0] data_ram_6_dina; // @[dcache.scala 111:65]
  wire [31:0] data_ram_6_douta; // @[dcache.scala 111:65]
  wire [3:0] data_ram_6_wea; // @[dcache.scala 111:65]
  wire [7:0] data_ram_7_addra; // @[dcache.scala 111:65]
  wire  data_ram_7_clka; // @[dcache.scala 111:65]
  wire [31:0] data_ram_7_dina; // @[dcache.scala 111:65]
  wire [31:0] data_ram_7_douta; // @[dcache.scala 111:65]
  wire [3:0] data_ram_7_wea; // @[dcache.scala 111:65]
  wire  LFSR_result_prng_clock; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_reset; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_5; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_6; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_7; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_8; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_9; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_10; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_11; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_12; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_13; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_14; // @[PRNG.scala 91:22]
  wire  LFSR_result_prng_io_out_15; // @[PRNG.scala 91:22]
  wire  _cacheOperation_T_1 = 3'h0 == cache_op; // @[Lookup.scala 31:38]
  wire  _cacheOperation_T_3 = 3'h1 == cache_op; // @[Lookup.scala 31:38]
  wire  _cacheOperation_T_5 = 3'h2 == cache_op; // @[Lookup.scala 31:38]
  wire  _cacheOperation_T_7 = 3'h3 == cache_op; // @[Lookup.scala 31:38]
  wire  _cacheOperation_T_9 = 3'h4 == cache_op; // @[Lookup.scala 31:38]
  wire  _cacheOperation_T_11 = 3'h5 == cache_op; // @[Lookup.scala 31:38]
  wire  _cacheOperation_T_13 = 3'h6 == cache_op; // @[Lookup.scala 31:38]
  wire  _cacheOperation_T_20 = _cacheOperation_T_7 ? 1'h0 : _cacheOperation_T_9 | _cacheOperation_T_11; // @[Lookup.scala 34:39]
  wire  _cacheOperation_T_21 = _cacheOperation_T_5 ? 1'h0 : _cacheOperation_T_20; // @[Lookup.scala 34:39]
  wire  _cacheOperation_T_22 = _cacheOperation_T_3 ? 1'h0 : _cacheOperation_T_21; // @[Lookup.scala 34:39]
  wire  cacheOperation_0 = _cacheOperation_T_1 | _cacheOperation_T_22; // @[Lookup.scala 34:39]
  wire  _cacheOperation_T_36 = _cacheOperation_T_3 ? 1'h0 : _cacheOperation_T_5; // @[Lookup.scala 34:39]
  wire  _cacheOperation_T_40 = _cacheOperation_T_9 ? 1'h0 : _cacheOperation_T_11 | _cacheOperation_T_13; // @[Lookup.scala 34:39]
  wire  _cacheOperation_T_41 = _cacheOperation_T_7 ? 1'h0 : _cacheOperation_T_40; // @[Lookup.scala 34:39]
  wire  _cacheOperation_T_42 = _cacheOperation_T_5 ? 1'h0 : _cacheOperation_T_41; // @[Lookup.scala 34:39]
  wire  _cacheOperation_T_43 = _cacheOperation_T_3 ? 1'h0 : _cacheOperation_T_42; // @[Lookup.scala 34:39]
  wire  cacheOperation_3 = _cacheOperation_T_1 | _cacheOperation_T_43; // @[Lookup.scala 34:39]
  wire  cacheOperation_4 = _cacheOperation_T_1 | (_cacheOperation_T_3 | _cacheOperation_T_5); // @[Lookup.scala 34:39]
  reg  cacheInst_r; // @[dcache.scala 89:38]
  reg  invalidate; // @[dcache.scala 90:38]
  reg  loadTag; // @[dcache.scala 91:38]
  reg  storeTag; // @[dcache.scala 92:38]
  reg  writeBack; // @[dcache.scala 93:38]
  reg  indexOnly; // @[dcache.scala 94:38]
  reg  dirty_0_0; // @[dcache.scala 113:28]
  reg  dirty_0_1; // @[dcache.scala 113:28]
  reg  dirty_0_2; // @[dcache.scala 113:28]
  reg  dirty_0_3; // @[dcache.scala 113:28]
  reg  dirty_0_4; // @[dcache.scala 113:28]
  reg  dirty_0_5; // @[dcache.scala 113:28]
  reg  dirty_0_6; // @[dcache.scala 113:28]
  reg  dirty_0_7; // @[dcache.scala 113:28]
  reg  dirty_0_8; // @[dcache.scala 113:28]
  reg  dirty_0_9; // @[dcache.scala 113:28]
  reg  dirty_0_10; // @[dcache.scala 113:28]
  reg  dirty_0_11; // @[dcache.scala 113:28]
  reg  dirty_0_12; // @[dcache.scala 113:28]
  reg  dirty_0_13; // @[dcache.scala 113:28]
  reg  dirty_0_14; // @[dcache.scala 113:28]
  reg  dirty_0_15; // @[dcache.scala 113:28]
  reg  dirty_0_16; // @[dcache.scala 113:28]
  reg  dirty_0_17; // @[dcache.scala 113:28]
  reg  dirty_0_18; // @[dcache.scala 113:28]
  reg  dirty_0_19; // @[dcache.scala 113:28]
  reg  dirty_0_20; // @[dcache.scala 113:28]
  reg  dirty_0_21; // @[dcache.scala 113:28]
  reg  dirty_0_22; // @[dcache.scala 113:28]
  reg  dirty_0_23; // @[dcache.scala 113:28]
  reg  dirty_0_24; // @[dcache.scala 113:28]
  reg  dirty_0_25; // @[dcache.scala 113:28]
  reg  dirty_0_26; // @[dcache.scala 113:28]
  reg  dirty_0_27; // @[dcache.scala 113:28]
  reg  dirty_0_28; // @[dcache.scala 113:28]
  reg  dirty_0_29; // @[dcache.scala 113:28]
  reg  dirty_0_30; // @[dcache.scala 113:28]
  reg  dirty_0_31; // @[dcache.scala 113:28]
  reg  dirty_0_32; // @[dcache.scala 113:28]
  reg  dirty_0_33; // @[dcache.scala 113:28]
  reg  dirty_0_34; // @[dcache.scala 113:28]
  reg  dirty_0_35; // @[dcache.scala 113:28]
  reg  dirty_0_36; // @[dcache.scala 113:28]
  reg  dirty_0_37; // @[dcache.scala 113:28]
  reg  dirty_0_38; // @[dcache.scala 113:28]
  reg  dirty_0_39; // @[dcache.scala 113:28]
  reg  dirty_0_40; // @[dcache.scala 113:28]
  reg  dirty_0_41; // @[dcache.scala 113:28]
  reg  dirty_0_42; // @[dcache.scala 113:28]
  reg  dirty_0_43; // @[dcache.scala 113:28]
  reg  dirty_0_44; // @[dcache.scala 113:28]
  reg  dirty_0_45; // @[dcache.scala 113:28]
  reg  dirty_0_46; // @[dcache.scala 113:28]
  reg  dirty_0_47; // @[dcache.scala 113:28]
  reg  dirty_0_48; // @[dcache.scala 113:28]
  reg  dirty_0_49; // @[dcache.scala 113:28]
  reg  dirty_0_50; // @[dcache.scala 113:28]
  reg  dirty_0_51; // @[dcache.scala 113:28]
  reg  dirty_0_52; // @[dcache.scala 113:28]
  reg  dirty_0_53; // @[dcache.scala 113:28]
  reg  dirty_0_54; // @[dcache.scala 113:28]
  reg  dirty_0_55; // @[dcache.scala 113:28]
  reg  dirty_0_56; // @[dcache.scala 113:28]
  reg  dirty_0_57; // @[dcache.scala 113:28]
  reg  dirty_0_58; // @[dcache.scala 113:28]
  reg  dirty_0_59; // @[dcache.scala 113:28]
  reg  dirty_0_60; // @[dcache.scala 113:28]
  reg  dirty_0_61; // @[dcache.scala 113:28]
  reg  dirty_0_62; // @[dcache.scala 113:28]
  reg  dirty_0_63; // @[dcache.scala 113:28]
  reg  dirty_0_64; // @[dcache.scala 113:28]
  reg  dirty_0_65; // @[dcache.scala 113:28]
  reg  dirty_0_66; // @[dcache.scala 113:28]
  reg  dirty_0_67; // @[dcache.scala 113:28]
  reg  dirty_0_68; // @[dcache.scala 113:28]
  reg  dirty_0_69; // @[dcache.scala 113:28]
  reg  dirty_0_70; // @[dcache.scala 113:28]
  reg  dirty_0_71; // @[dcache.scala 113:28]
  reg  dirty_0_72; // @[dcache.scala 113:28]
  reg  dirty_0_73; // @[dcache.scala 113:28]
  reg  dirty_0_74; // @[dcache.scala 113:28]
  reg  dirty_0_75; // @[dcache.scala 113:28]
  reg  dirty_0_76; // @[dcache.scala 113:28]
  reg  dirty_0_77; // @[dcache.scala 113:28]
  reg  dirty_0_78; // @[dcache.scala 113:28]
  reg  dirty_0_79; // @[dcache.scala 113:28]
  reg  dirty_0_80; // @[dcache.scala 113:28]
  reg  dirty_0_81; // @[dcache.scala 113:28]
  reg  dirty_0_82; // @[dcache.scala 113:28]
  reg  dirty_0_83; // @[dcache.scala 113:28]
  reg  dirty_0_84; // @[dcache.scala 113:28]
  reg  dirty_0_85; // @[dcache.scala 113:28]
  reg  dirty_0_86; // @[dcache.scala 113:28]
  reg  dirty_0_87; // @[dcache.scala 113:28]
  reg  dirty_0_88; // @[dcache.scala 113:28]
  reg  dirty_0_89; // @[dcache.scala 113:28]
  reg  dirty_0_90; // @[dcache.scala 113:28]
  reg  dirty_0_91; // @[dcache.scala 113:28]
  reg  dirty_0_92; // @[dcache.scala 113:28]
  reg  dirty_0_93; // @[dcache.scala 113:28]
  reg  dirty_0_94; // @[dcache.scala 113:28]
  reg  dirty_0_95; // @[dcache.scala 113:28]
  reg  dirty_0_96; // @[dcache.scala 113:28]
  reg  dirty_0_97; // @[dcache.scala 113:28]
  reg  dirty_0_98; // @[dcache.scala 113:28]
  reg  dirty_0_99; // @[dcache.scala 113:28]
  reg  dirty_0_100; // @[dcache.scala 113:28]
  reg  dirty_0_101; // @[dcache.scala 113:28]
  reg  dirty_0_102; // @[dcache.scala 113:28]
  reg  dirty_0_103; // @[dcache.scala 113:28]
  reg  dirty_0_104; // @[dcache.scala 113:28]
  reg  dirty_0_105; // @[dcache.scala 113:28]
  reg  dirty_0_106; // @[dcache.scala 113:28]
  reg  dirty_0_107; // @[dcache.scala 113:28]
  reg  dirty_0_108; // @[dcache.scala 113:28]
  reg  dirty_0_109; // @[dcache.scala 113:28]
  reg  dirty_0_110; // @[dcache.scala 113:28]
  reg  dirty_0_111; // @[dcache.scala 113:28]
  reg  dirty_0_112; // @[dcache.scala 113:28]
  reg  dirty_0_113; // @[dcache.scala 113:28]
  reg  dirty_0_114; // @[dcache.scala 113:28]
  reg  dirty_0_115; // @[dcache.scala 113:28]
  reg  dirty_0_116; // @[dcache.scala 113:28]
  reg  dirty_0_117; // @[dcache.scala 113:28]
  reg  dirty_0_118; // @[dcache.scala 113:28]
  reg  dirty_0_119; // @[dcache.scala 113:28]
  reg  dirty_0_120; // @[dcache.scala 113:28]
  reg  dirty_0_121; // @[dcache.scala 113:28]
  reg  dirty_0_122; // @[dcache.scala 113:28]
  reg  dirty_0_123; // @[dcache.scala 113:28]
  reg  dirty_0_124; // @[dcache.scala 113:28]
  reg  dirty_0_125; // @[dcache.scala 113:28]
  reg  dirty_0_126; // @[dcache.scala 113:28]
  reg  dirty_0_127; // @[dcache.scala 113:28]
  reg  dirty_0_128; // @[dcache.scala 113:28]
  reg  dirty_0_129; // @[dcache.scala 113:28]
  reg  dirty_0_130; // @[dcache.scala 113:28]
  reg  dirty_0_131; // @[dcache.scala 113:28]
  reg  dirty_0_132; // @[dcache.scala 113:28]
  reg  dirty_0_133; // @[dcache.scala 113:28]
  reg  dirty_0_134; // @[dcache.scala 113:28]
  reg  dirty_0_135; // @[dcache.scala 113:28]
  reg  dirty_0_136; // @[dcache.scala 113:28]
  reg  dirty_0_137; // @[dcache.scala 113:28]
  reg  dirty_0_138; // @[dcache.scala 113:28]
  reg  dirty_0_139; // @[dcache.scala 113:28]
  reg  dirty_0_140; // @[dcache.scala 113:28]
  reg  dirty_0_141; // @[dcache.scala 113:28]
  reg  dirty_0_142; // @[dcache.scala 113:28]
  reg  dirty_0_143; // @[dcache.scala 113:28]
  reg  dirty_0_144; // @[dcache.scala 113:28]
  reg  dirty_0_145; // @[dcache.scala 113:28]
  reg  dirty_0_146; // @[dcache.scala 113:28]
  reg  dirty_0_147; // @[dcache.scala 113:28]
  reg  dirty_0_148; // @[dcache.scala 113:28]
  reg  dirty_0_149; // @[dcache.scala 113:28]
  reg  dirty_0_150; // @[dcache.scala 113:28]
  reg  dirty_0_151; // @[dcache.scala 113:28]
  reg  dirty_0_152; // @[dcache.scala 113:28]
  reg  dirty_0_153; // @[dcache.scala 113:28]
  reg  dirty_0_154; // @[dcache.scala 113:28]
  reg  dirty_0_155; // @[dcache.scala 113:28]
  reg  dirty_0_156; // @[dcache.scala 113:28]
  reg  dirty_0_157; // @[dcache.scala 113:28]
  reg  dirty_0_158; // @[dcache.scala 113:28]
  reg  dirty_0_159; // @[dcache.scala 113:28]
  reg  dirty_0_160; // @[dcache.scala 113:28]
  reg  dirty_0_161; // @[dcache.scala 113:28]
  reg  dirty_0_162; // @[dcache.scala 113:28]
  reg  dirty_0_163; // @[dcache.scala 113:28]
  reg  dirty_0_164; // @[dcache.scala 113:28]
  reg  dirty_0_165; // @[dcache.scala 113:28]
  reg  dirty_0_166; // @[dcache.scala 113:28]
  reg  dirty_0_167; // @[dcache.scala 113:28]
  reg  dirty_0_168; // @[dcache.scala 113:28]
  reg  dirty_0_169; // @[dcache.scala 113:28]
  reg  dirty_0_170; // @[dcache.scala 113:28]
  reg  dirty_0_171; // @[dcache.scala 113:28]
  reg  dirty_0_172; // @[dcache.scala 113:28]
  reg  dirty_0_173; // @[dcache.scala 113:28]
  reg  dirty_0_174; // @[dcache.scala 113:28]
  reg  dirty_0_175; // @[dcache.scala 113:28]
  reg  dirty_0_176; // @[dcache.scala 113:28]
  reg  dirty_0_177; // @[dcache.scala 113:28]
  reg  dirty_0_178; // @[dcache.scala 113:28]
  reg  dirty_0_179; // @[dcache.scala 113:28]
  reg  dirty_0_180; // @[dcache.scala 113:28]
  reg  dirty_0_181; // @[dcache.scala 113:28]
  reg  dirty_0_182; // @[dcache.scala 113:28]
  reg  dirty_0_183; // @[dcache.scala 113:28]
  reg  dirty_0_184; // @[dcache.scala 113:28]
  reg  dirty_0_185; // @[dcache.scala 113:28]
  reg  dirty_0_186; // @[dcache.scala 113:28]
  reg  dirty_0_187; // @[dcache.scala 113:28]
  reg  dirty_0_188; // @[dcache.scala 113:28]
  reg  dirty_0_189; // @[dcache.scala 113:28]
  reg  dirty_0_190; // @[dcache.scala 113:28]
  reg  dirty_0_191; // @[dcache.scala 113:28]
  reg  dirty_0_192; // @[dcache.scala 113:28]
  reg  dirty_0_193; // @[dcache.scala 113:28]
  reg  dirty_0_194; // @[dcache.scala 113:28]
  reg  dirty_0_195; // @[dcache.scala 113:28]
  reg  dirty_0_196; // @[dcache.scala 113:28]
  reg  dirty_0_197; // @[dcache.scala 113:28]
  reg  dirty_0_198; // @[dcache.scala 113:28]
  reg  dirty_0_199; // @[dcache.scala 113:28]
  reg  dirty_0_200; // @[dcache.scala 113:28]
  reg  dirty_0_201; // @[dcache.scala 113:28]
  reg  dirty_0_202; // @[dcache.scala 113:28]
  reg  dirty_0_203; // @[dcache.scala 113:28]
  reg  dirty_0_204; // @[dcache.scala 113:28]
  reg  dirty_0_205; // @[dcache.scala 113:28]
  reg  dirty_0_206; // @[dcache.scala 113:28]
  reg  dirty_0_207; // @[dcache.scala 113:28]
  reg  dirty_0_208; // @[dcache.scala 113:28]
  reg  dirty_0_209; // @[dcache.scala 113:28]
  reg  dirty_0_210; // @[dcache.scala 113:28]
  reg  dirty_0_211; // @[dcache.scala 113:28]
  reg  dirty_0_212; // @[dcache.scala 113:28]
  reg  dirty_0_213; // @[dcache.scala 113:28]
  reg  dirty_0_214; // @[dcache.scala 113:28]
  reg  dirty_0_215; // @[dcache.scala 113:28]
  reg  dirty_0_216; // @[dcache.scala 113:28]
  reg  dirty_0_217; // @[dcache.scala 113:28]
  reg  dirty_0_218; // @[dcache.scala 113:28]
  reg  dirty_0_219; // @[dcache.scala 113:28]
  reg  dirty_0_220; // @[dcache.scala 113:28]
  reg  dirty_0_221; // @[dcache.scala 113:28]
  reg  dirty_0_222; // @[dcache.scala 113:28]
  reg  dirty_0_223; // @[dcache.scala 113:28]
  reg  dirty_0_224; // @[dcache.scala 113:28]
  reg  dirty_0_225; // @[dcache.scala 113:28]
  reg  dirty_0_226; // @[dcache.scala 113:28]
  reg  dirty_0_227; // @[dcache.scala 113:28]
  reg  dirty_0_228; // @[dcache.scala 113:28]
  reg  dirty_0_229; // @[dcache.scala 113:28]
  reg  dirty_0_230; // @[dcache.scala 113:28]
  reg  dirty_0_231; // @[dcache.scala 113:28]
  reg  dirty_0_232; // @[dcache.scala 113:28]
  reg  dirty_0_233; // @[dcache.scala 113:28]
  reg  dirty_0_234; // @[dcache.scala 113:28]
  reg  dirty_0_235; // @[dcache.scala 113:28]
  reg  dirty_0_236; // @[dcache.scala 113:28]
  reg  dirty_0_237; // @[dcache.scala 113:28]
  reg  dirty_0_238; // @[dcache.scala 113:28]
  reg  dirty_0_239; // @[dcache.scala 113:28]
  reg  dirty_0_240; // @[dcache.scala 113:28]
  reg  dirty_0_241; // @[dcache.scala 113:28]
  reg  dirty_0_242; // @[dcache.scala 113:28]
  reg  dirty_0_243; // @[dcache.scala 113:28]
  reg  dirty_0_244; // @[dcache.scala 113:28]
  reg  dirty_0_245; // @[dcache.scala 113:28]
  reg  dirty_0_246; // @[dcache.scala 113:28]
  reg  dirty_0_247; // @[dcache.scala 113:28]
  reg  dirty_0_248; // @[dcache.scala 113:28]
  reg  dirty_0_249; // @[dcache.scala 113:28]
  reg  dirty_0_250; // @[dcache.scala 113:28]
  reg  dirty_0_251; // @[dcache.scala 113:28]
  reg  dirty_0_252; // @[dcache.scala 113:28]
  reg  dirty_0_253; // @[dcache.scala 113:28]
  reg  dirty_0_254; // @[dcache.scala 113:28]
  reg  dirty_0_255; // @[dcache.scala 113:28]
  reg  dirty_1_0; // @[dcache.scala 113:28]
  reg  dirty_1_1; // @[dcache.scala 113:28]
  reg  dirty_1_2; // @[dcache.scala 113:28]
  reg  dirty_1_3; // @[dcache.scala 113:28]
  reg  dirty_1_4; // @[dcache.scala 113:28]
  reg  dirty_1_5; // @[dcache.scala 113:28]
  reg  dirty_1_6; // @[dcache.scala 113:28]
  reg  dirty_1_7; // @[dcache.scala 113:28]
  reg  dirty_1_8; // @[dcache.scala 113:28]
  reg  dirty_1_9; // @[dcache.scala 113:28]
  reg  dirty_1_10; // @[dcache.scala 113:28]
  reg  dirty_1_11; // @[dcache.scala 113:28]
  reg  dirty_1_12; // @[dcache.scala 113:28]
  reg  dirty_1_13; // @[dcache.scala 113:28]
  reg  dirty_1_14; // @[dcache.scala 113:28]
  reg  dirty_1_15; // @[dcache.scala 113:28]
  reg  dirty_1_16; // @[dcache.scala 113:28]
  reg  dirty_1_17; // @[dcache.scala 113:28]
  reg  dirty_1_18; // @[dcache.scala 113:28]
  reg  dirty_1_19; // @[dcache.scala 113:28]
  reg  dirty_1_20; // @[dcache.scala 113:28]
  reg  dirty_1_21; // @[dcache.scala 113:28]
  reg  dirty_1_22; // @[dcache.scala 113:28]
  reg  dirty_1_23; // @[dcache.scala 113:28]
  reg  dirty_1_24; // @[dcache.scala 113:28]
  reg  dirty_1_25; // @[dcache.scala 113:28]
  reg  dirty_1_26; // @[dcache.scala 113:28]
  reg  dirty_1_27; // @[dcache.scala 113:28]
  reg  dirty_1_28; // @[dcache.scala 113:28]
  reg  dirty_1_29; // @[dcache.scala 113:28]
  reg  dirty_1_30; // @[dcache.scala 113:28]
  reg  dirty_1_31; // @[dcache.scala 113:28]
  reg  dirty_1_32; // @[dcache.scala 113:28]
  reg  dirty_1_33; // @[dcache.scala 113:28]
  reg  dirty_1_34; // @[dcache.scala 113:28]
  reg  dirty_1_35; // @[dcache.scala 113:28]
  reg  dirty_1_36; // @[dcache.scala 113:28]
  reg  dirty_1_37; // @[dcache.scala 113:28]
  reg  dirty_1_38; // @[dcache.scala 113:28]
  reg  dirty_1_39; // @[dcache.scala 113:28]
  reg  dirty_1_40; // @[dcache.scala 113:28]
  reg  dirty_1_41; // @[dcache.scala 113:28]
  reg  dirty_1_42; // @[dcache.scala 113:28]
  reg  dirty_1_43; // @[dcache.scala 113:28]
  reg  dirty_1_44; // @[dcache.scala 113:28]
  reg  dirty_1_45; // @[dcache.scala 113:28]
  reg  dirty_1_46; // @[dcache.scala 113:28]
  reg  dirty_1_47; // @[dcache.scala 113:28]
  reg  dirty_1_48; // @[dcache.scala 113:28]
  reg  dirty_1_49; // @[dcache.scala 113:28]
  reg  dirty_1_50; // @[dcache.scala 113:28]
  reg  dirty_1_51; // @[dcache.scala 113:28]
  reg  dirty_1_52; // @[dcache.scala 113:28]
  reg  dirty_1_53; // @[dcache.scala 113:28]
  reg  dirty_1_54; // @[dcache.scala 113:28]
  reg  dirty_1_55; // @[dcache.scala 113:28]
  reg  dirty_1_56; // @[dcache.scala 113:28]
  reg  dirty_1_57; // @[dcache.scala 113:28]
  reg  dirty_1_58; // @[dcache.scala 113:28]
  reg  dirty_1_59; // @[dcache.scala 113:28]
  reg  dirty_1_60; // @[dcache.scala 113:28]
  reg  dirty_1_61; // @[dcache.scala 113:28]
  reg  dirty_1_62; // @[dcache.scala 113:28]
  reg  dirty_1_63; // @[dcache.scala 113:28]
  reg  dirty_1_64; // @[dcache.scala 113:28]
  reg  dirty_1_65; // @[dcache.scala 113:28]
  reg  dirty_1_66; // @[dcache.scala 113:28]
  reg  dirty_1_67; // @[dcache.scala 113:28]
  reg  dirty_1_68; // @[dcache.scala 113:28]
  reg  dirty_1_69; // @[dcache.scala 113:28]
  reg  dirty_1_70; // @[dcache.scala 113:28]
  reg  dirty_1_71; // @[dcache.scala 113:28]
  reg  dirty_1_72; // @[dcache.scala 113:28]
  reg  dirty_1_73; // @[dcache.scala 113:28]
  reg  dirty_1_74; // @[dcache.scala 113:28]
  reg  dirty_1_75; // @[dcache.scala 113:28]
  reg  dirty_1_76; // @[dcache.scala 113:28]
  reg  dirty_1_77; // @[dcache.scala 113:28]
  reg  dirty_1_78; // @[dcache.scala 113:28]
  reg  dirty_1_79; // @[dcache.scala 113:28]
  reg  dirty_1_80; // @[dcache.scala 113:28]
  reg  dirty_1_81; // @[dcache.scala 113:28]
  reg  dirty_1_82; // @[dcache.scala 113:28]
  reg  dirty_1_83; // @[dcache.scala 113:28]
  reg  dirty_1_84; // @[dcache.scala 113:28]
  reg  dirty_1_85; // @[dcache.scala 113:28]
  reg  dirty_1_86; // @[dcache.scala 113:28]
  reg  dirty_1_87; // @[dcache.scala 113:28]
  reg  dirty_1_88; // @[dcache.scala 113:28]
  reg  dirty_1_89; // @[dcache.scala 113:28]
  reg  dirty_1_90; // @[dcache.scala 113:28]
  reg  dirty_1_91; // @[dcache.scala 113:28]
  reg  dirty_1_92; // @[dcache.scala 113:28]
  reg  dirty_1_93; // @[dcache.scala 113:28]
  reg  dirty_1_94; // @[dcache.scala 113:28]
  reg  dirty_1_95; // @[dcache.scala 113:28]
  reg  dirty_1_96; // @[dcache.scala 113:28]
  reg  dirty_1_97; // @[dcache.scala 113:28]
  reg  dirty_1_98; // @[dcache.scala 113:28]
  reg  dirty_1_99; // @[dcache.scala 113:28]
  reg  dirty_1_100; // @[dcache.scala 113:28]
  reg  dirty_1_101; // @[dcache.scala 113:28]
  reg  dirty_1_102; // @[dcache.scala 113:28]
  reg  dirty_1_103; // @[dcache.scala 113:28]
  reg  dirty_1_104; // @[dcache.scala 113:28]
  reg  dirty_1_105; // @[dcache.scala 113:28]
  reg  dirty_1_106; // @[dcache.scala 113:28]
  reg  dirty_1_107; // @[dcache.scala 113:28]
  reg  dirty_1_108; // @[dcache.scala 113:28]
  reg  dirty_1_109; // @[dcache.scala 113:28]
  reg  dirty_1_110; // @[dcache.scala 113:28]
  reg  dirty_1_111; // @[dcache.scala 113:28]
  reg  dirty_1_112; // @[dcache.scala 113:28]
  reg  dirty_1_113; // @[dcache.scala 113:28]
  reg  dirty_1_114; // @[dcache.scala 113:28]
  reg  dirty_1_115; // @[dcache.scala 113:28]
  reg  dirty_1_116; // @[dcache.scala 113:28]
  reg  dirty_1_117; // @[dcache.scala 113:28]
  reg  dirty_1_118; // @[dcache.scala 113:28]
  reg  dirty_1_119; // @[dcache.scala 113:28]
  reg  dirty_1_120; // @[dcache.scala 113:28]
  reg  dirty_1_121; // @[dcache.scala 113:28]
  reg  dirty_1_122; // @[dcache.scala 113:28]
  reg  dirty_1_123; // @[dcache.scala 113:28]
  reg  dirty_1_124; // @[dcache.scala 113:28]
  reg  dirty_1_125; // @[dcache.scala 113:28]
  reg  dirty_1_126; // @[dcache.scala 113:28]
  reg  dirty_1_127; // @[dcache.scala 113:28]
  reg  dirty_1_128; // @[dcache.scala 113:28]
  reg  dirty_1_129; // @[dcache.scala 113:28]
  reg  dirty_1_130; // @[dcache.scala 113:28]
  reg  dirty_1_131; // @[dcache.scala 113:28]
  reg  dirty_1_132; // @[dcache.scala 113:28]
  reg  dirty_1_133; // @[dcache.scala 113:28]
  reg  dirty_1_134; // @[dcache.scala 113:28]
  reg  dirty_1_135; // @[dcache.scala 113:28]
  reg  dirty_1_136; // @[dcache.scala 113:28]
  reg  dirty_1_137; // @[dcache.scala 113:28]
  reg  dirty_1_138; // @[dcache.scala 113:28]
  reg  dirty_1_139; // @[dcache.scala 113:28]
  reg  dirty_1_140; // @[dcache.scala 113:28]
  reg  dirty_1_141; // @[dcache.scala 113:28]
  reg  dirty_1_142; // @[dcache.scala 113:28]
  reg  dirty_1_143; // @[dcache.scala 113:28]
  reg  dirty_1_144; // @[dcache.scala 113:28]
  reg  dirty_1_145; // @[dcache.scala 113:28]
  reg  dirty_1_146; // @[dcache.scala 113:28]
  reg  dirty_1_147; // @[dcache.scala 113:28]
  reg  dirty_1_148; // @[dcache.scala 113:28]
  reg  dirty_1_149; // @[dcache.scala 113:28]
  reg  dirty_1_150; // @[dcache.scala 113:28]
  reg  dirty_1_151; // @[dcache.scala 113:28]
  reg  dirty_1_152; // @[dcache.scala 113:28]
  reg  dirty_1_153; // @[dcache.scala 113:28]
  reg  dirty_1_154; // @[dcache.scala 113:28]
  reg  dirty_1_155; // @[dcache.scala 113:28]
  reg  dirty_1_156; // @[dcache.scala 113:28]
  reg  dirty_1_157; // @[dcache.scala 113:28]
  reg  dirty_1_158; // @[dcache.scala 113:28]
  reg  dirty_1_159; // @[dcache.scala 113:28]
  reg  dirty_1_160; // @[dcache.scala 113:28]
  reg  dirty_1_161; // @[dcache.scala 113:28]
  reg  dirty_1_162; // @[dcache.scala 113:28]
  reg  dirty_1_163; // @[dcache.scala 113:28]
  reg  dirty_1_164; // @[dcache.scala 113:28]
  reg  dirty_1_165; // @[dcache.scala 113:28]
  reg  dirty_1_166; // @[dcache.scala 113:28]
  reg  dirty_1_167; // @[dcache.scala 113:28]
  reg  dirty_1_168; // @[dcache.scala 113:28]
  reg  dirty_1_169; // @[dcache.scala 113:28]
  reg  dirty_1_170; // @[dcache.scala 113:28]
  reg  dirty_1_171; // @[dcache.scala 113:28]
  reg  dirty_1_172; // @[dcache.scala 113:28]
  reg  dirty_1_173; // @[dcache.scala 113:28]
  reg  dirty_1_174; // @[dcache.scala 113:28]
  reg  dirty_1_175; // @[dcache.scala 113:28]
  reg  dirty_1_176; // @[dcache.scala 113:28]
  reg  dirty_1_177; // @[dcache.scala 113:28]
  reg  dirty_1_178; // @[dcache.scala 113:28]
  reg  dirty_1_179; // @[dcache.scala 113:28]
  reg  dirty_1_180; // @[dcache.scala 113:28]
  reg  dirty_1_181; // @[dcache.scala 113:28]
  reg  dirty_1_182; // @[dcache.scala 113:28]
  reg  dirty_1_183; // @[dcache.scala 113:28]
  reg  dirty_1_184; // @[dcache.scala 113:28]
  reg  dirty_1_185; // @[dcache.scala 113:28]
  reg  dirty_1_186; // @[dcache.scala 113:28]
  reg  dirty_1_187; // @[dcache.scala 113:28]
  reg  dirty_1_188; // @[dcache.scala 113:28]
  reg  dirty_1_189; // @[dcache.scala 113:28]
  reg  dirty_1_190; // @[dcache.scala 113:28]
  reg  dirty_1_191; // @[dcache.scala 113:28]
  reg  dirty_1_192; // @[dcache.scala 113:28]
  reg  dirty_1_193; // @[dcache.scala 113:28]
  reg  dirty_1_194; // @[dcache.scala 113:28]
  reg  dirty_1_195; // @[dcache.scala 113:28]
  reg  dirty_1_196; // @[dcache.scala 113:28]
  reg  dirty_1_197; // @[dcache.scala 113:28]
  reg  dirty_1_198; // @[dcache.scala 113:28]
  reg  dirty_1_199; // @[dcache.scala 113:28]
  reg  dirty_1_200; // @[dcache.scala 113:28]
  reg  dirty_1_201; // @[dcache.scala 113:28]
  reg  dirty_1_202; // @[dcache.scala 113:28]
  reg  dirty_1_203; // @[dcache.scala 113:28]
  reg  dirty_1_204; // @[dcache.scala 113:28]
  reg  dirty_1_205; // @[dcache.scala 113:28]
  reg  dirty_1_206; // @[dcache.scala 113:28]
  reg  dirty_1_207; // @[dcache.scala 113:28]
  reg  dirty_1_208; // @[dcache.scala 113:28]
  reg  dirty_1_209; // @[dcache.scala 113:28]
  reg  dirty_1_210; // @[dcache.scala 113:28]
  reg  dirty_1_211; // @[dcache.scala 113:28]
  reg  dirty_1_212; // @[dcache.scala 113:28]
  reg  dirty_1_213; // @[dcache.scala 113:28]
  reg  dirty_1_214; // @[dcache.scala 113:28]
  reg  dirty_1_215; // @[dcache.scala 113:28]
  reg  dirty_1_216; // @[dcache.scala 113:28]
  reg  dirty_1_217; // @[dcache.scala 113:28]
  reg  dirty_1_218; // @[dcache.scala 113:28]
  reg  dirty_1_219; // @[dcache.scala 113:28]
  reg  dirty_1_220; // @[dcache.scala 113:28]
  reg  dirty_1_221; // @[dcache.scala 113:28]
  reg  dirty_1_222; // @[dcache.scala 113:28]
  reg  dirty_1_223; // @[dcache.scala 113:28]
  reg  dirty_1_224; // @[dcache.scala 113:28]
  reg  dirty_1_225; // @[dcache.scala 113:28]
  reg  dirty_1_226; // @[dcache.scala 113:28]
  reg  dirty_1_227; // @[dcache.scala 113:28]
  reg  dirty_1_228; // @[dcache.scala 113:28]
  reg  dirty_1_229; // @[dcache.scala 113:28]
  reg  dirty_1_230; // @[dcache.scala 113:28]
  reg  dirty_1_231; // @[dcache.scala 113:28]
  reg  dirty_1_232; // @[dcache.scala 113:28]
  reg  dirty_1_233; // @[dcache.scala 113:28]
  reg  dirty_1_234; // @[dcache.scala 113:28]
  reg  dirty_1_235; // @[dcache.scala 113:28]
  reg  dirty_1_236; // @[dcache.scala 113:28]
  reg  dirty_1_237; // @[dcache.scala 113:28]
  reg  dirty_1_238; // @[dcache.scala 113:28]
  reg  dirty_1_239; // @[dcache.scala 113:28]
  reg  dirty_1_240; // @[dcache.scala 113:28]
  reg  dirty_1_241; // @[dcache.scala 113:28]
  reg  dirty_1_242; // @[dcache.scala 113:28]
  reg  dirty_1_243; // @[dcache.scala 113:28]
  reg  dirty_1_244; // @[dcache.scala 113:28]
  reg  dirty_1_245; // @[dcache.scala 113:28]
  reg  dirty_1_246; // @[dcache.scala 113:28]
  reg  dirty_1_247; // @[dcache.scala 113:28]
  reg  dirty_1_248; // @[dcache.scala 113:28]
  reg  dirty_1_249; // @[dcache.scala 113:28]
  reg  dirty_1_250; // @[dcache.scala 113:28]
  reg  dirty_1_251; // @[dcache.scala 113:28]
  reg  dirty_1_252; // @[dcache.scala 113:28]
  reg  dirty_1_253; // @[dcache.scala 113:28]
  reg  dirty_1_254; // @[dcache.scala 113:28]
  reg  dirty_1_255; // @[dcache.scala 113:28]
  reg  req_valid; // @[dcache.scala 116:34]
  reg  req_op; // @[dcache.scala 118:34]
  reg  req_uncached; // @[dcache.scala 119:34]
  reg [3:0] req_offset; // @[dcache.scala 120:34]
  reg [2:0] req_lstype; // @[dcache.scala 121:34]
  reg [7:0] req_set; // @[dcache.scala 122:34]
  reg [19:0] req_tag; // @[dcache.scala 123:34]
  reg [3:0] req_wstrb_0; // @[dcache.scala 124:34]
  reg [31:0] req_wdata_0; // @[dcache.scala 125:34]
  reg [31:0] req_wdata_1; // @[dcache.scala 127:34]
  reg [3:0] req_wstrb_1; // @[dcache.scala 128:34]
  reg  req_wline; // @[dcache.scala 129:34]
  reg [7:0] req_wset; // @[dcache.scala 130:34]
  reg [3:0] req_woffset; // @[dcache.scala 131:34]
  reg [20:0] tagv_r_0; // @[dcache.scala 136:34]
  reg [20:0] tagv_r_1; // @[dcache.scala 136:34]
  wire  waySel = req_tag[0]; // @[dcache.scala 137:31]
  reg [2:0] state; // @[dcache.scala 171:34]
  reg  refillIDX_r; // @[dcache.scala 174:34]
  wire [7:0] LFSR_result_lo = {LFSR_result_prng_io_out_7,LFSR_result_prng_io_out_6,LFSR_result_prng_io_out_5,
    LFSR_result_prng_io_out_4,LFSR_result_prng_io_out_3,LFSR_result_prng_io_out_2,LFSR_result_prng_io_out_1,
    LFSR_result_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [7:0] LFSR_result_hi = {LFSR_result_prng_io_out_15,LFSR_result_prng_io_out_14,LFSR_result_prng_io_out_13,
    LFSR_result_prng_io_out_12,LFSR_result_prng_io_out_11,LFSR_result_prng_io_out_10,LFSR_result_prng_io_out_9,
    LFSR_result_prng_io_out_8}; // @[PRNG.scala 95:17]
  reg [15:0] LFSR_result; // @[dcache.scala 177:34]
  reg [1:0] wr_cnt; // @[dcache.scala 178:34]
  wire [2:0] _state_T = uncached ? 3'h3 : 3'h1; // @[dcache.scala 205:39]
  wire  _GEN_2 = valid ? op : req_op; // @[dcache.scala 204:30 207:33 118:34]
  wire [19:0] _GEN_4 = valid ? tag : req_tag; // @[dcache.scala 204:30 209:33 123:34]
  wire [7:0] _GEN_5 = valid ? index : req_set; // @[dcache.scala 204:30 210:33 122:34]
  wire [3:0] _GEN_6 = valid ? offset : req_offset; // @[dcache.scala 204:30 211:33 120:34]
  wire  _GEN_7 = valid ? uncached : req_uncached; // @[dcache.scala 204:30 212:33 119:34]
  wire [2:0] _GEN_8 = valid ? lstype : req_lstype; // @[dcache.scala 204:30 213:33 121:34]
  wire [3:0] _GEN_9 = valid ? wstrb : req_wstrb_0; // @[dcache.scala 204:30 214:33 124:34]
  wire [31:0] _GEN_10 = valid ? wdata : req_wdata_0; // @[dcache.scala 204:30 215:33 125:34]
  wire [7:0] _GEN_15 = cache_op_en ? cache_index : _GEN_5; // @[dcache.scala 185:30 190:33]
  wire  _GEN_22 = cache_op_en ? 1'h0 : valid; // @[dcache.scala 156:25 185:30]
  wire [20:0] tagv_0_douta = tagv_ram_douta; // @[dcache.scala 110:{42,42}]
  wire  _hit_T = ~req_uncached; // @[dcache.scala 227:36]
  wire [31:0] data_0_0_douta = data_ram_douta; // @[dcache.scala 111:{58,58}]
  wire [31:0] data_0_1_douta = data_ram_1_douta; // @[dcache.scala 111:{58,58}]
  wire [31:0] _GEN_29 = 2'h1 == req_offset[3:2] ? data_0_1_douta : data_0_0_douta; // @[dcache.scala 228:{33,33}]
  wire [31:0] data_0_2_douta = data_ram_2_douta; // @[dcache.scala 111:{58,58}]
  wire [31:0] _GEN_30 = 2'h2 == req_offset[3:2] ? data_0_2_douta : _GEN_29; // @[dcache.scala 228:{33,33}]
  wire [31:0] data_0_3_douta = data_ram_3_douta; // @[dcache.scala 111:{58,58}]
  wire [31:0] _GEN_31 = 2'h3 == req_offset[3:2] ? data_0_3_douta : _GEN_30; // @[dcache.scala 228:{33,33}]
  wire  _T_6 = ~req_op; // @[dcache.scala 229:26]
  wire  _T_7 = ~cacheInst_r; // @[dcache.scala 233:31]
  wire [3:0] _GEN_32 = ~cacheInst_r ? req_offset : req_woffset; // @[dcache.scala 131:34 233:44 234:37]
  wire [7:0] _GEN_33 = ~cacheInst_r ? req_set : req_wset; // @[dcache.scala 130:34 233:44 235:37]
  wire  _GEN_34 = ~cacheInst_r ? 1'h0 : req_wline; // @[dcache.scala 129:34 233:44 236:37]
  wire [3:0] _GEN_35 = ~cacheInst_r ? req_wstrb_0 : req_wstrb_1; // @[dcache.scala 128:34 233:44 237:37]
  wire [31:0] _GEN_36 = ~cacheInst_r ? req_wdata_0 : req_wdata_1; // @[dcache.scala 127:34 233:44 238:37]
  wire [3:0] _GEN_38 = _T_6 ? req_woffset : _GEN_32; // @[dcache.scala 230:21 131:34]
  wire [7:0] _GEN_39 = _T_6 ? req_wset : _GEN_33; // @[dcache.scala 230:21 130:34]
  wire  _GEN_40 = _T_6 ? req_wline : _GEN_34; // @[dcache.scala 230:21 129:34]
  wire [3:0] _GEN_41 = _T_6 ? req_wstrb_1 : _GEN_35; // @[dcache.scala 230:21 128:34]
  wire [31:0] _GEN_42 = _T_6 ? req_wdata_1 : _GEN_36; // @[dcache.scala 230:21 127:34]
  wire  _GEN_43 = ~indexOnly ? 1'h0 : refillIDX_r; // @[dcache.scala 174:34 240:37 241:37]
  reg [1:0] wstate; // @[dcache.scala 441:31]
  wire [20:0] tagv_1_douta = tagv_ram_1_douta; // @[dcache.scala 110:{42,42}]
  wire  _GEN_74 = tagv_1_douta[19:0] == req_tag & tagv_1_douta[20] & _T_6; // @[dcache.scala 226:78]
  wire  _GEN_8082 = 3'h3 == state & refillIDX_r; // @[dcache.scala 183:18 335:23 167:25]
  wire  _GEN_8639 = 3'h2 == state ? 1'h0 : _GEN_8082; // @[dcache.scala 183:18 167:25]
  wire  _GEN_9194 = 3'h1 == state ? _GEN_74 : _GEN_8639; // @[dcache.scala 183:18]
  wire  req_rline = 3'h0 == state ? 1'h0 : _GEN_9194; // @[dcache.scala 183:18 167:25]
  reg  req_wline_1; // @[dcache.scala 444:32]
  reg [3:0] req_woffset_1; // @[dcache.scala 443:32]
  wire  _war_stall_T_22 = _T_6 & state == 3'h1 & (req_woffset[3:2] == req_offset[3:2] | req_woffset_1[3:2] == req_offset
    [3:2]) | state == 3'h2; // @[dcache.scala 477:127]
  wire  war_stall = (wstate == 2'h1 | wstate == 2'h2) & req_valid & _hit_T & (req_wline == req_rline | req_wline_1 ==
    req_rline) & _war_stall_T_22; // @[dcache.scala 476:165]
  wire  _T_9 = ~war_stall; // @[dcache.scala 244:26]
  wire  _T_11 = ~war_stall & _T_7; // @[dcache.scala 244:37]
  wire  _GEN_45 = tagv_0_douta[19:0] == req_tag & tagv_0_douta[20] & ~req_uncached; // @[dcache.scala 154:25 226:78 227:33]
  wire [31:0] _GEN_46 = tagv_0_douta[19:0] == req_tag & tagv_0_douta[20] ? _GEN_31 : 32'h7777; // @[dcache.scala 155:25 226:78 228:33]
  wire [3:0] _GEN_48 = tagv_0_douta[19:0] == req_tag & tagv_0_douta[20] ? _GEN_38 : req_woffset; // @[dcache.scala 131:34 226:78]
  wire [7:0] _GEN_49 = tagv_0_douta[19:0] == req_tag & tagv_0_douta[20] ? _GEN_39 : req_wset; // @[dcache.scala 130:34 226:78]
  wire  _GEN_50 = tagv_0_douta[19:0] == req_tag & tagv_0_douta[20] ? _GEN_40 : req_wline; // @[dcache.scala 129:34 226:78]
  wire [3:0] _GEN_51 = tagv_0_douta[19:0] == req_tag & tagv_0_douta[20] ? _GEN_41 : req_wstrb_1; // @[dcache.scala 128:34 226:78]
  wire [31:0] _GEN_52 = tagv_0_douta[19:0] == req_tag & tagv_0_douta[20] ? _GEN_42 : req_wdata_1; // @[dcache.scala 127:34 226:78]
  wire  _GEN_53 = tagv_0_douta[19:0] == req_tag & tagv_0_douta[20] ? _GEN_43 : refillIDX_r; // @[dcache.scala 174:34 226:78]
  wire  _GEN_54 = tagv_0_douta[19:0] == req_tag & tagv_0_douta[20] & _T_11; // @[dcache.scala 157:25 226:78]
  wire [31:0] data_1_0_douta = data_ram_4_douta; // @[dcache.scala 111:{58,58}]
  wire [31:0] data_1_1_douta = data_ram_5_douta; // @[dcache.scala 111:{58,58}]
  wire [31:0] _GEN_56 = 2'h1 == req_offset[3:2] ? data_1_1_douta : data_1_0_douta; // @[dcache.scala 228:{33,33}]
  wire [31:0] data_1_2_douta = data_ram_6_douta; // @[dcache.scala 111:{58,58}]
  wire [31:0] _GEN_57 = 2'h2 == req_offset[3:2] ? data_1_2_douta : _GEN_56; // @[dcache.scala 228:{33,33}]
  wire [31:0] data_1_3_douta = data_ram_7_douta; // @[dcache.scala 111:{58,58}]
  wire [31:0] _GEN_58 = 2'h3 == req_offset[3:2] ? data_1_3_douta : _GEN_57; // @[dcache.scala 228:{33,33}]
  wire [3:0] _GEN_59 = ~cacheInst_r ? req_offset : _GEN_48; // @[dcache.scala 233:44 234:37]
  wire [7:0] _GEN_60 = ~cacheInst_r ? req_set : _GEN_49; // @[dcache.scala 233:44 235:37]
  wire  _GEN_61 = ~cacheInst_r | _GEN_50; // @[dcache.scala 233:44 236:37]
  wire [3:0] _GEN_62 = ~cacheInst_r ? req_wstrb_0 : _GEN_51; // @[dcache.scala 233:44 237:37]
  wire [31:0] _GEN_63 = ~cacheInst_r ? req_wdata_0 : _GEN_52; // @[dcache.scala 233:44 238:37]
  wire [3:0] _GEN_65 = _T_6 ? _GEN_48 : _GEN_59; // @[dcache.scala 230:21]
  wire [7:0] _GEN_66 = _T_6 ? _GEN_49 : _GEN_60; // @[dcache.scala 230:21]
  wire  _GEN_67 = _T_6 ? _GEN_50 : _GEN_61; // @[dcache.scala 230:21]
  wire [3:0] _GEN_68 = _T_6 ? _GEN_51 : _GEN_62; // @[dcache.scala 230:21]
  wire [31:0] _GEN_69 = _T_6 ? _GEN_52 : _GEN_63; // @[dcache.scala 230:21]
  wire  _GEN_70 = ~indexOnly | _GEN_53; // @[dcache.scala 240:37 241:37]
  wire  _GEN_71 = _T_11 | _GEN_54; // @[dcache.scala 245:21 246:37]
  wire  _GEN_72 = tagv_1_douta[19:0] == req_tag & tagv_1_douta[20] ? ~req_uncached : _GEN_45; // @[dcache.scala 226:78 227:33]
  wire [31:0] _GEN_73 = tagv_1_douta[19:0] == req_tag & tagv_1_douta[20] ? _GEN_58 : _GEN_46; // @[dcache.scala 226:78 228:33]
  wire  _GEN_80 = tagv_1_douta[19:0] == req_tag & tagv_1_douta[20] ? _GEN_70 : _GEN_53; // @[dcache.scala 226:78]
  wire  _GEN_81 = tagv_1_douta[19:0] == req_tag & tagv_1_douta[20] ? _GEN_71 : _GEN_54; // @[dcache.scala 226:78]
  wire [2:0] _state_T_1 = storeTag ? 3'h5 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _state_T_2 = loadTag ? 3'h5 : _state_T_1; // @[Mux.scala 101:16]
  wire [2:0] _state_T_3 = invalidate ? 3'h5 : _state_T_2; // @[Mux.scala 101:16]
  wire [2:0] _state_T_4 = writeBack ? 3'h3 : _state_T_3; // @[Mux.scala 101:16]
  wire [2:0] _state_T_5 = invalidate ? 3'h5 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _state_T_6 = writeBack ? 3'h3 : _state_T_5; // @[Mux.scala 101:16]
  wire [2:0] _GEN_82 = hit ? _state_T_6 : 3'h0; // @[dcache.scala 265:31 266:33 279:37]
  wire  _GEN_83 = hit ? 1'h0 : 1'h1; // @[dcache.scala 265:31 97:21 272:37]
  wire  _GEN_84 = hit & cacheInst_r; // @[dcache.scala 265:31 273:37 89:38]
  wire  _GEN_85 = hit & invalidate; // @[dcache.scala 265:31 274:37 90:38]
  wire  _GEN_86 = hit & indexOnly; // @[dcache.scala 265:31 275:37 94:38]
  wire  _GEN_87 = hit & writeBack; // @[dcache.scala 265:31 276:37 93:38]
  wire  _GEN_88 = hit & storeTag; // @[dcache.scala 265:31 277:37 92:38]
  wire  _GEN_89 = hit & loadTag; // @[dcache.scala 265:31 278:37 91:38]
  wire [2:0] _GEN_90 = indexOnly ? _state_T_4 : _GEN_82; // @[dcache.scala 256:32 257:33]
  wire  _GEN_91 = indexOnly ? waySel : _GEN_80; // @[dcache.scala 256:32 263:37]
  wire  _GEN_92 = indexOnly ? 1'h0 : _GEN_83; // @[dcache.scala 256:32 97:21]
  wire  _GEN_93 = indexOnly ? cacheInst_r : _GEN_84; // @[dcache.scala 256:32 89:38]
  wire  _GEN_94 = indexOnly ? invalidate : _GEN_85; // @[dcache.scala 256:32 90:38]
  wire  _GEN_95 = indexOnly ? indexOnly : _GEN_86; // @[dcache.scala 256:32 94:38]
  wire  _GEN_96 = indexOnly ? writeBack : _GEN_87; // @[dcache.scala 256:32 93:38]
  wire  _GEN_97 = indexOnly ? storeTag : _GEN_88; // @[dcache.scala 256:32 92:38]
  wire  _GEN_98 = indexOnly ? loadTag : _GEN_89; // @[dcache.scala 256:32 91:38]
  wire [2:0] _GEN_99 = valid ? _state_T : 3'h0; // @[dcache.scala 287:19 288:39 307:29]
  wire [2:0] _GEN_101 = _T_9 ? _GEN_99 : 3'h1; // @[dcache.scala 285:34 311:27]
  wire  _GEN_102 = _T_9 & valid; // @[dcache.scala 156:25 285:34]
  wire  _GEN_103 = _T_9 ? valid : req_valid; // @[dcache.scala 116:34 285:34]
  wire  _GEN_104 = _T_9 ? _GEN_7 : req_uncached; // @[dcache.scala 119:34 285:34]
  wire [2:0] _GEN_105 = _T_9 ? _GEN_8 : req_lstype; // @[dcache.scala 121:34 285:34]
  wire  _GEN_106 = _T_9 ? _GEN_2 : req_op; // @[dcache.scala 118:34 285:34]
  wire [19:0] _GEN_107 = _T_9 ? _GEN_4 : req_tag; // @[dcache.scala 123:34 285:34]
  wire [7:0] _GEN_108 = _T_9 ? _GEN_5 : req_set; // @[dcache.scala 122:34 285:34]
  wire [3:0] _GEN_109 = _T_9 ? _GEN_6 : req_offset; // @[dcache.scala 120:34 285:34]
  wire [3:0] _GEN_110 = _T_9 ? _GEN_9 : req_wstrb_0; // @[dcache.scala 124:34 285:34]
  wire [31:0] _GEN_111 = _T_9 ? _GEN_10 : req_wdata_0; // @[dcache.scala 125:34 285:34]
  wire [2:0] _GEN_112 = ~hit ? 3'h2 : _GEN_101; // @[dcache.scala 282:28 283:33]
  wire  _GEN_113 = ~hit ? 1'h0 : _GEN_102; // @[dcache.scala 156:25 282:28]
  wire  _GEN_114 = ~hit ? req_valid : _GEN_103; // @[dcache.scala 282:28 116:34]
  wire  _GEN_115 = ~hit ? req_uncached : _GEN_104; // @[dcache.scala 282:28 119:34]
  wire [2:0] _GEN_116 = ~hit ? req_lstype : _GEN_105; // @[dcache.scala 282:28 121:34]
  wire  _GEN_117 = ~hit ? req_op : _GEN_106; // @[dcache.scala 282:28 118:34]
  wire [19:0] _GEN_118 = ~hit ? req_tag : _GEN_107; // @[dcache.scala 282:28 123:34]
  wire [7:0] _GEN_119 = ~hit ? req_set : _GEN_108; // @[dcache.scala 282:28 122:34]
  wire [3:0] _GEN_120 = ~hit ? req_offset : _GEN_109; // @[dcache.scala 282:28 120:34]
  wire [3:0] _GEN_121 = ~hit ? req_wstrb_0 : _GEN_110; // @[dcache.scala 282:28 124:34]
  wire [31:0] _GEN_122 = ~hit ? req_wdata_0 : _GEN_111; // @[dcache.scala 282:28 125:34]
  wire  _GEN_125 = cacheInst_r & _GEN_92; // @[dcache.scala 255:30 97:21]
  wire  _GEN_132 = cacheInst_r ? 1'h0 : _GEN_113; // @[dcache.scala 156:25 255:30]
  wire [7:0] _GEN_138 = cacheInst_r ? req_set : _GEN_119; // @[dcache.scala 255:30 122:34]
  wire  _T_28 = ~tagv_r_1[20]; // @[dcache.scala 317:22]
  wire  _GEN_144 = ~tagv_r_1[20] | ~tagv_r_0[20]; // @[dcache.scala 317:37 318:41]
  wire  _GEN_147 = tagv_r_0[19:0] == req_tag & tagv_r_0[20] ? 1'h0 : _T_28; // @[dcache.scala 323:68 325:41]
  wire  _GEN_148 = tagv_r_1[19:0] == req_tag & tagv_r_1[20] | (tagv_r_0[19:0] == req_tag & tagv_r_0[20] | _GEN_144); // @[dcache.scala 323:68 324:41]
  wire  _GEN_149 = tagv_r_1[19:0] == req_tag & tagv_r_1[20] | _GEN_147; // @[dcache.scala 323:68 325:41]
  wire  _GEN_9222 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_148; // @[dcache.scala 183:18 180:25]
  wire  refillHit = 3'h0 == state ? 1'h0 : _GEN_9222; // @[dcache.scala 183:18 180:25]
  wire  _GEN_150 = ~refillHit ? LFSR_result[0] : _GEN_149; // @[dcache.scala 328:30 329:27]
  wire  _GEN_11958 = ~refillIDX_r; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11959 = 8'h1 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_152 = ~refillIDX_r & 8'h1 == req_set ? dirty_0_1 : dirty_0_0; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11961 = 8'h2 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_153 = ~refillIDX_r & 8'h2 == req_set ? dirty_0_2 : _GEN_152; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11963 = 8'h3 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_154 = ~refillIDX_r & 8'h3 == req_set ? dirty_0_3 : _GEN_153; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11965 = 8'h4 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_155 = ~refillIDX_r & 8'h4 == req_set ? dirty_0_4 : _GEN_154; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11967 = 8'h5 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_156 = ~refillIDX_r & 8'h5 == req_set ? dirty_0_5 : _GEN_155; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11969 = 8'h6 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_157 = ~refillIDX_r & 8'h6 == req_set ? dirty_0_6 : _GEN_156; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11971 = 8'h7 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_158 = ~refillIDX_r & 8'h7 == req_set ? dirty_0_7 : _GEN_157; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11973 = 8'h8 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_159 = ~refillIDX_r & 8'h8 == req_set ? dirty_0_8 : _GEN_158; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11975 = 8'h9 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_160 = ~refillIDX_r & 8'h9 == req_set ? dirty_0_9 : _GEN_159; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11977 = 8'ha == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_161 = ~refillIDX_r & 8'ha == req_set ? dirty_0_10 : _GEN_160; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11979 = 8'hb == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_162 = ~refillIDX_r & 8'hb == req_set ? dirty_0_11 : _GEN_161; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11981 = 8'hc == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_163 = ~refillIDX_r & 8'hc == req_set ? dirty_0_12 : _GEN_162; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11983 = 8'hd == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_164 = ~refillIDX_r & 8'hd == req_set ? dirty_0_13 : _GEN_163; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11985 = 8'he == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_165 = ~refillIDX_r & 8'he == req_set ? dirty_0_14 : _GEN_164; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11987 = 8'hf == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_166 = ~refillIDX_r & 8'hf == req_set ? dirty_0_15 : _GEN_165; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11989 = 8'h10 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_167 = ~refillIDX_r & 8'h10 == req_set ? dirty_0_16 : _GEN_166; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11991 = 8'h11 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_168 = ~refillIDX_r & 8'h11 == req_set ? dirty_0_17 : _GEN_167; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11993 = 8'h12 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_169 = ~refillIDX_r & 8'h12 == req_set ? dirty_0_18 : _GEN_168; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11995 = 8'h13 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_170 = ~refillIDX_r & 8'h13 == req_set ? dirty_0_19 : _GEN_169; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11997 = 8'h14 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_171 = ~refillIDX_r & 8'h14 == req_set ? dirty_0_20 : _GEN_170; // @[dcache.scala 345:{54,54}]
  wire  _GEN_11999 = 8'h15 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_172 = ~refillIDX_r & 8'h15 == req_set ? dirty_0_21 : _GEN_171; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12001 = 8'h16 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_173 = ~refillIDX_r & 8'h16 == req_set ? dirty_0_22 : _GEN_172; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12003 = 8'h17 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_174 = ~refillIDX_r & 8'h17 == req_set ? dirty_0_23 : _GEN_173; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12005 = 8'h18 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_175 = ~refillIDX_r & 8'h18 == req_set ? dirty_0_24 : _GEN_174; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12007 = 8'h19 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_176 = ~refillIDX_r & 8'h19 == req_set ? dirty_0_25 : _GEN_175; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12009 = 8'h1a == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_177 = ~refillIDX_r & 8'h1a == req_set ? dirty_0_26 : _GEN_176; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12011 = 8'h1b == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_178 = ~refillIDX_r & 8'h1b == req_set ? dirty_0_27 : _GEN_177; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12013 = 8'h1c == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_179 = ~refillIDX_r & 8'h1c == req_set ? dirty_0_28 : _GEN_178; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12015 = 8'h1d == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_180 = ~refillIDX_r & 8'h1d == req_set ? dirty_0_29 : _GEN_179; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12017 = 8'h1e == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_181 = ~refillIDX_r & 8'h1e == req_set ? dirty_0_30 : _GEN_180; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12019 = 8'h1f == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_182 = ~refillIDX_r & 8'h1f == req_set ? dirty_0_31 : _GEN_181; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12021 = 8'h20 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_183 = ~refillIDX_r & 8'h20 == req_set ? dirty_0_32 : _GEN_182; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12023 = 8'h21 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_184 = ~refillIDX_r & 8'h21 == req_set ? dirty_0_33 : _GEN_183; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12025 = 8'h22 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_185 = ~refillIDX_r & 8'h22 == req_set ? dirty_0_34 : _GEN_184; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12027 = 8'h23 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_186 = ~refillIDX_r & 8'h23 == req_set ? dirty_0_35 : _GEN_185; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12029 = 8'h24 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_187 = ~refillIDX_r & 8'h24 == req_set ? dirty_0_36 : _GEN_186; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12031 = 8'h25 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_188 = ~refillIDX_r & 8'h25 == req_set ? dirty_0_37 : _GEN_187; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12033 = 8'h26 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_189 = ~refillIDX_r & 8'h26 == req_set ? dirty_0_38 : _GEN_188; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12035 = 8'h27 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_190 = ~refillIDX_r & 8'h27 == req_set ? dirty_0_39 : _GEN_189; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12037 = 8'h28 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_191 = ~refillIDX_r & 8'h28 == req_set ? dirty_0_40 : _GEN_190; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12039 = 8'h29 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_192 = ~refillIDX_r & 8'h29 == req_set ? dirty_0_41 : _GEN_191; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12041 = 8'h2a == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_193 = ~refillIDX_r & 8'h2a == req_set ? dirty_0_42 : _GEN_192; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12043 = 8'h2b == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_194 = ~refillIDX_r & 8'h2b == req_set ? dirty_0_43 : _GEN_193; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12045 = 8'h2c == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_195 = ~refillIDX_r & 8'h2c == req_set ? dirty_0_44 : _GEN_194; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12047 = 8'h2d == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_196 = ~refillIDX_r & 8'h2d == req_set ? dirty_0_45 : _GEN_195; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12049 = 8'h2e == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_197 = ~refillIDX_r & 8'h2e == req_set ? dirty_0_46 : _GEN_196; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12051 = 8'h2f == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_198 = ~refillIDX_r & 8'h2f == req_set ? dirty_0_47 : _GEN_197; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12053 = 8'h30 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_199 = ~refillIDX_r & 8'h30 == req_set ? dirty_0_48 : _GEN_198; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12055 = 8'h31 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_200 = ~refillIDX_r & 8'h31 == req_set ? dirty_0_49 : _GEN_199; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12057 = 8'h32 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_201 = ~refillIDX_r & 8'h32 == req_set ? dirty_0_50 : _GEN_200; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12059 = 8'h33 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_202 = ~refillIDX_r & 8'h33 == req_set ? dirty_0_51 : _GEN_201; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12061 = 8'h34 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_203 = ~refillIDX_r & 8'h34 == req_set ? dirty_0_52 : _GEN_202; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12063 = 8'h35 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_204 = ~refillIDX_r & 8'h35 == req_set ? dirty_0_53 : _GEN_203; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12065 = 8'h36 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_205 = ~refillIDX_r & 8'h36 == req_set ? dirty_0_54 : _GEN_204; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12067 = 8'h37 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_206 = ~refillIDX_r & 8'h37 == req_set ? dirty_0_55 : _GEN_205; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12069 = 8'h38 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_207 = ~refillIDX_r & 8'h38 == req_set ? dirty_0_56 : _GEN_206; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12071 = 8'h39 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_208 = ~refillIDX_r & 8'h39 == req_set ? dirty_0_57 : _GEN_207; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12073 = 8'h3a == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_209 = ~refillIDX_r & 8'h3a == req_set ? dirty_0_58 : _GEN_208; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12075 = 8'h3b == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_210 = ~refillIDX_r & 8'h3b == req_set ? dirty_0_59 : _GEN_209; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12077 = 8'h3c == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_211 = ~refillIDX_r & 8'h3c == req_set ? dirty_0_60 : _GEN_210; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12079 = 8'h3d == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_212 = ~refillIDX_r & 8'h3d == req_set ? dirty_0_61 : _GEN_211; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12081 = 8'h3e == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_213 = ~refillIDX_r & 8'h3e == req_set ? dirty_0_62 : _GEN_212; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12083 = 8'h3f == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_214 = ~refillIDX_r & 8'h3f == req_set ? dirty_0_63 : _GEN_213; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12085 = 8'h40 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_215 = ~refillIDX_r & 8'h40 == req_set ? dirty_0_64 : _GEN_214; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12087 = 8'h41 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_216 = ~refillIDX_r & 8'h41 == req_set ? dirty_0_65 : _GEN_215; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12089 = 8'h42 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_217 = ~refillIDX_r & 8'h42 == req_set ? dirty_0_66 : _GEN_216; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12091 = 8'h43 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_218 = ~refillIDX_r & 8'h43 == req_set ? dirty_0_67 : _GEN_217; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12093 = 8'h44 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_219 = ~refillIDX_r & 8'h44 == req_set ? dirty_0_68 : _GEN_218; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12095 = 8'h45 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_220 = ~refillIDX_r & 8'h45 == req_set ? dirty_0_69 : _GEN_219; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12097 = 8'h46 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_221 = ~refillIDX_r & 8'h46 == req_set ? dirty_0_70 : _GEN_220; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12099 = 8'h47 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_222 = ~refillIDX_r & 8'h47 == req_set ? dirty_0_71 : _GEN_221; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12101 = 8'h48 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_223 = ~refillIDX_r & 8'h48 == req_set ? dirty_0_72 : _GEN_222; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12103 = 8'h49 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_224 = ~refillIDX_r & 8'h49 == req_set ? dirty_0_73 : _GEN_223; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12105 = 8'h4a == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_225 = ~refillIDX_r & 8'h4a == req_set ? dirty_0_74 : _GEN_224; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12107 = 8'h4b == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_226 = ~refillIDX_r & 8'h4b == req_set ? dirty_0_75 : _GEN_225; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12109 = 8'h4c == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_227 = ~refillIDX_r & 8'h4c == req_set ? dirty_0_76 : _GEN_226; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12111 = 8'h4d == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_228 = ~refillIDX_r & 8'h4d == req_set ? dirty_0_77 : _GEN_227; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12113 = 8'h4e == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_229 = ~refillIDX_r & 8'h4e == req_set ? dirty_0_78 : _GEN_228; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12115 = 8'h4f == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_230 = ~refillIDX_r & 8'h4f == req_set ? dirty_0_79 : _GEN_229; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12117 = 8'h50 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_231 = ~refillIDX_r & 8'h50 == req_set ? dirty_0_80 : _GEN_230; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12119 = 8'h51 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_232 = ~refillIDX_r & 8'h51 == req_set ? dirty_0_81 : _GEN_231; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12121 = 8'h52 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_233 = ~refillIDX_r & 8'h52 == req_set ? dirty_0_82 : _GEN_232; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12123 = 8'h53 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_234 = ~refillIDX_r & 8'h53 == req_set ? dirty_0_83 : _GEN_233; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12125 = 8'h54 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_235 = ~refillIDX_r & 8'h54 == req_set ? dirty_0_84 : _GEN_234; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12127 = 8'h55 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_236 = ~refillIDX_r & 8'h55 == req_set ? dirty_0_85 : _GEN_235; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12129 = 8'h56 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_237 = ~refillIDX_r & 8'h56 == req_set ? dirty_0_86 : _GEN_236; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12131 = 8'h57 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_238 = ~refillIDX_r & 8'h57 == req_set ? dirty_0_87 : _GEN_237; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12133 = 8'h58 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_239 = ~refillIDX_r & 8'h58 == req_set ? dirty_0_88 : _GEN_238; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12135 = 8'h59 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_240 = ~refillIDX_r & 8'h59 == req_set ? dirty_0_89 : _GEN_239; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12137 = 8'h5a == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_241 = ~refillIDX_r & 8'h5a == req_set ? dirty_0_90 : _GEN_240; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12139 = 8'h5b == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_242 = ~refillIDX_r & 8'h5b == req_set ? dirty_0_91 : _GEN_241; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12141 = 8'h5c == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_243 = ~refillIDX_r & 8'h5c == req_set ? dirty_0_92 : _GEN_242; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12143 = 8'h5d == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_244 = ~refillIDX_r & 8'h5d == req_set ? dirty_0_93 : _GEN_243; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12145 = 8'h5e == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_245 = ~refillIDX_r & 8'h5e == req_set ? dirty_0_94 : _GEN_244; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12147 = 8'h5f == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_246 = ~refillIDX_r & 8'h5f == req_set ? dirty_0_95 : _GEN_245; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12149 = 8'h60 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_247 = ~refillIDX_r & 8'h60 == req_set ? dirty_0_96 : _GEN_246; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12151 = 8'h61 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_248 = ~refillIDX_r & 8'h61 == req_set ? dirty_0_97 : _GEN_247; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12153 = 8'h62 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_249 = ~refillIDX_r & 8'h62 == req_set ? dirty_0_98 : _GEN_248; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12155 = 8'h63 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_250 = ~refillIDX_r & 8'h63 == req_set ? dirty_0_99 : _GEN_249; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12157 = 8'h64 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_251 = ~refillIDX_r & 8'h64 == req_set ? dirty_0_100 : _GEN_250; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12159 = 8'h65 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_252 = ~refillIDX_r & 8'h65 == req_set ? dirty_0_101 : _GEN_251; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12161 = 8'h66 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_253 = ~refillIDX_r & 8'h66 == req_set ? dirty_0_102 : _GEN_252; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12163 = 8'h67 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_254 = ~refillIDX_r & 8'h67 == req_set ? dirty_0_103 : _GEN_253; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12165 = 8'h68 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_255 = ~refillIDX_r & 8'h68 == req_set ? dirty_0_104 : _GEN_254; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12167 = 8'h69 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_256 = ~refillIDX_r & 8'h69 == req_set ? dirty_0_105 : _GEN_255; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12169 = 8'h6a == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_257 = ~refillIDX_r & 8'h6a == req_set ? dirty_0_106 : _GEN_256; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12171 = 8'h6b == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_258 = ~refillIDX_r & 8'h6b == req_set ? dirty_0_107 : _GEN_257; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12173 = 8'h6c == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_259 = ~refillIDX_r & 8'h6c == req_set ? dirty_0_108 : _GEN_258; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12175 = 8'h6d == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_260 = ~refillIDX_r & 8'h6d == req_set ? dirty_0_109 : _GEN_259; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12177 = 8'h6e == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_261 = ~refillIDX_r & 8'h6e == req_set ? dirty_0_110 : _GEN_260; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12179 = 8'h6f == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_262 = ~refillIDX_r & 8'h6f == req_set ? dirty_0_111 : _GEN_261; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12181 = 8'h70 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_263 = ~refillIDX_r & 8'h70 == req_set ? dirty_0_112 : _GEN_262; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12183 = 8'h71 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_264 = ~refillIDX_r & 8'h71 == req_set ? dirty_0_113 : _GEN_263; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12185 = 8'h72 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_265 = ~refillIDX_r & 8'h72 == req_set ? dirty_0_114 : _GEN_264; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12187 = 8'h73 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_266 = ~refillIDX_r & 8'h73 == req_set ? dirty_0_115 : _GEN_265; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12189 = 8'h74 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_267 = ~refillIDX_r & 8'h74 == req_set ? dirty_0_116 : _GEN_266; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12191 = 8'h75 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_268 = ~refillIDX_r & 8'h75 == req_set ? dirty_0_117 : _GEN_267; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12193 = 8'h76 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_269 = ~refillIDX_r & 8'h76 == req_set ? dirty_0_118 : _GEN_268; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12195 = 8'h77 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_270 = ~refillIDX_r & 8'h77 == req_set ? dirty_0_119 : _GEN_269; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12197 = 8'h78 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_271 = ~refillIDX_r & 8'h78 == req_set ? dirty_0_120 : _GEN_270; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12199 = 8'h79 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_272 = ~refillIDX_r & 8'h79 == req_set ? dirty_0_121 : _GEN_271; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12201 = 8'h7a == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_273 = ~refillIDX_r & 8'h7a == req_set ? dirty_0_122 : _GEN_272; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12203 = 8'h7b == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_274 = ~refillIDX_r & 8'h7b == req_set ? dirty_0_123 : _GEN_273; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12205 = 8'h7c == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_275 = ~refillIDX_r & 8'h7c == req_set ? dirty_0_124 : _GEN_274; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12207 = 8'h7d == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_276 = ~refillIDX_r & 8'h7d == req_set ? dirty_0_125 : _GEN_275; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12209 = 8'h7e == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_277 = ~refillIDX_r & 8'h7e == req_set ? dirty_0_126 : _GEN_276; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12211 = 8'h7f == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_278 = ~refillIDX_r & 8'h7f == req_set ? dirty_0_127 : _GEN_277; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12213 = 8'h80 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_279 = ~refillIDX_r & 8'h80 == req_set ? dirty_0_128 : _GEN_278; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12215 = 8'h81 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_280 = ~refillIDX_r & 8'h81 == req_set ? dirty_0_129 : _GEN_279; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12217 = 8'h82 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_281 = ~refillIDX_r & 8'h82 == req_set ? dirty_0_130 : _GEN_280; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12219 = 8'h83 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_282 = ~refillIDX_r & 8'h83 == req_set ? dirty_0_131 : _GEN_281; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12221 = 8'h84 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_283 = ~refillIDX_r & 8'h84 == req_set ? dirty_0_132 : _GEN_282; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12223 = 8'h85 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_284 = ~refillIDX_r & 8'h85 == req_set ? dirty_0_133 : _GEN_283; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12225 = 8'h86 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_285 = ~refillIDX_r & 8'h86 == req_set ? dirty_0_134 : _GEN_284; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12227 = 8'h87 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_286 = ~refillIDX_r & 8'h87 == req_set ? dirty_0_135 : _GEN_285; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12229 = 8'h88 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_287 = ~refillIDX_r & 8'h88 == req_set ? dirty_0_136 : _GEN_286; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12231 = 8'h89 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_288 = ~refillIDX_r & 8'h89 == req_set ? dirty_0_137 : _GEN_287; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12233 = 8'h8a == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_289 = ~refillIDX_r & 8'h8a == req_set ? dirty_0_138 : _GEN_288; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12235 = 8'h8b == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_290 = ~refillIDX_r & 8'h8b == req_set ? dirty_0_139 : _GEN_289; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12237 = 8'h8c == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_291 = ~refillIDX_r & 8'h8c == req_set ? dirty_0_140 : _GEN_290; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12239 = 8'h8d == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_292 = ~refillIDX_r & 8'h8d == req_set ? dirty_0_141 : _GEN_291; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12241 = 8'h8e == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_293 = ~refillIDX_r & 8'h8e == req_set ? dirty_0_142 : _GEN_292; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12243 = 8'h8f == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_294 = ~refillIDX_r & 8'h8f == req_set ? dirty_0_143 : _GEN_293; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12245 = 8'h90 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_295 = ~refillIDX_r & 8'h90 == req_set ? dirty_0_144 : _GEN_294; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12247 = 8'h91 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_296 = ~refillIDX_r & 8'h91 == req_set ? dirty_0_145 : _GEN_295; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12249 = 8'h92 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_297 = ~refillIDX_r & 8'h92 == req_set ? dirty_0_146 : _GEN_296; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12251 = 8'h93 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_298 = ~refillIDX_r & 8'h93 == req_set ? dirty_0_147 : _GEN_297; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12253 = 8'h94 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_299 = ~refillIDX_r & 8'h94 == req_set ? dirty_0_148 : _GEN_298; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12255 = 8'h95 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_300 = ~refillIDX_r & 8'h95 == req_set ? dirty_0_149 : _GEN_299; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12257 = 8'h96 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_301 = ~refillIDX_r & 8'h96 == req_set ? dirty_0_150 : _GEN_300; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12259 = 8'h97 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_302 = ~refillIDX_r & 8'h97 == req_set ? dirty_0_151 : _GEN_301; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12261 = 8'h98 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_303 = ~refillIDX_r & 8'h98 == req_set ? dirty_0_152 : _GEN_302; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12263 = 8'h99 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_304 = ~refillIDX_r & 8'h99 == req_set ? dirty_0_153 : _GEN_303; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12265 = 8'h9a == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_305 = ~refillIDX_r & 8'h9a == req_set ? dirty_0_154 : _GEN_304; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12267 = 8'h9b == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_306 = ~refillIDX_r & 8'h9b == req_set ? dirty_0_155 : _GEN_305; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12269 = 8'h9c == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_307 = ~refillIDX_r & 8'h9c == req_set ? dirty_0_156 : _GEN_306; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12271 = 8'h9d == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_308 = ~refillIDX_r & 8'h9d == req_set ? dirty_0_157 : _GEN_307; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12273 = 8'h9e == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_309 = ~refillIDX_r & 8'h9e == req_set ? dirty_0_158 : _GEN_308; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12275 = 8'h9f == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_310 = ~refillIDX_r & 8'h9f == req_set ? dirty_0_159 : _GEN_309; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12277 = 8'ha0 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_311 = ~refillIDX_r & 8'ha0 == req_set ? dirty_0_160 : _GEN_310; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12279 = 8'ha1 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_312 = ~refillIDX_r & 8'ha1 == req_set ? dirty_0_161 : _GEN_311; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12281 = 8'ha2 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_313 = ~refillIDX_r & 8'ha2 == req_set ? dirty_0_162 : _GEN_312; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12283 = 8'ha3 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_314 = ~refillIDX_r & 8'ha3 == req_set ? dirty_0_163 : _GEN_313; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12285 = 8'ha4 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_315 = ~refillIDX_r & 8'ha4 == req_set ? dirty_0_164 : _GEN_314; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12287 = 8'ha5 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_316 = ~refillIDX_r & 8'ha5 == req_set ? dirty_0_165 : _GEN_315; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12289 = 8'ha6 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_317 = ~refillIDX_r & 8'ha6 == req_set ? dirty_0_166 : _GEN_316; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12291 = 8'ha7 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_318 = ~refillIDX_r & 8'ha7 == req_set ? dirty_0_167 : _GEN_317; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12293 = 8'ha8 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_319 = ~refillIDX_r & 8'ha8 == req_set ? dirty_0_168 : _GEN_318; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12295 = 8'ha9 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_320 = ~refillIDX_r & 8'ha9 == req_set ? dirty_0_169 : _GEN_319; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12297 = 8'haa == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_321 = ~refillIDX_r & 8'haa == req_set ? dirty_0_170 : _GEN_320; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12299 = 8'hab == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_322 = ~refillIDX_r & 8'hab == req_set ? dirty_0_171 : _GEN_321; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12301 = 8'hac == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_323 = ~refillIDX_r & 8'hac == req_set ? dirty_0_172 : _GEN_322; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12303 = 8'had == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_324 = ~refillIDX_r & 8'had == req_set ? dirty_0_173 : _GEN_323; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12305 = 8'hae == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_325 = ~refillIDX_r & 8'hae == req_set ? dirty_0_174 : _GEN_324; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12307 = 8'haf == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_326 = ~refillIDX_r & 8'haf == req_set ? dirty_0_175 : _GEN_325; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12309 = 8'hb0 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_327 = ~refillIDX_r & 8'hb0 == req_set ? dirty_0_176 : _GEN_326; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12311 = 8'hb1 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_328 = ~refillIDX_r & 8'hb1 == req_set ? dirty_0_177 : _GEN_327; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12313 = 8'hb2 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_329 = ~refillIDX_r & 8'hb2 == req_set ? dirty_0_178 : _GEN_328; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12315 = 8'hb3 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_330 = ~refillIDX_r & 8'hb3 == req_set ? dirty_0_179 : _GEN_329; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12317 = 8'hb4 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_331 = ~refillIDX_r & 8'hb4 == req_set ? dirty_0_180 : _GEN_330; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12319 = 8'hb5 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_332 = ~refillIDX_r & 8'hb5 == req_set ? dirty_0_181 : _GEN_331; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12321 = 8'hb6 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_333 = ~refillIDX_r & 8'hb6 == req_set ? dirty_0_182 : _GEN_332; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12323 = 8'hb7 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_334 = ~refillIDX_r & 8'hb7 == req_set ? dirty_0_183 : _GEN_333; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12325 = 8'hb8 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_335 = ~refillIDX_r & 8'hb8 == req_set ? dirty_0_184 : _GEN_334; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12327 = 8'hb9 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_336 = ~refillIDX_r & 8'hb9 == req_set ? dirty_0_185 : _GEN_335; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12329 = 8'hba == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_337 = ~refillIDX_r & 8'hba == req_set ? dirty_0_186 : _GEN_336; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12331 = 8'hbb == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_338 = ~refillIDX_r & 8'hbb == req_set ? dirty_0_187 : _GEN_337; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12333 = 8'hbc == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_339 = ~refillIDX_r & 8'hbc == req_set ? dirty_0_188 : _GEN_338; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12335 = 8'hbd == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_340 = ~refillIDX_r & 8'hbd == req_set ? dirty_0_189 : _GEN_339; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12337 = 8'hbe == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_341 = ~refillIDX_r & 8'hbe == req_set ? dirty_0_190 : _GEN_340; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12339 = 8'hbf == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_342 = ~refillIDX_r & 8'hbf == req_set ? dirty_0_191 : _GEN_341; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12341 = 8'hc0 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_343 = ~refillIDX_r & 8'hc0 == req_set ? dirty_0_192 : _GEN_342; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12343 = 8'hc1 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_344 = ~refillIDX_r & 8'hc1 == req_set ? dirty_0_193 : _GEN_343; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12345 = 8'hc2 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_345 = ~refillIDX_r & 8'hc2 == req_set ? dirty_0_194 : _GEN_344; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12347 = 8'hc3 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_346 = ~refillIDX_r & 8'hc3 == req_set ? dirty_0_195 : _GEN_345; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12349 = 8'hc4 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_347 = ~refillIDX_r & 8'hc4 == req_set ? dirty_0_196 : _GEN_346; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12351 = 8'hc5 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_348 = ~refillIDX_r & 8'hc5 == req_set ? dirty_0_197 : _GEN_347; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12353 = 8'hc6 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_349 = ~refillIDX_r & 8'hc6 == req_set ? dirty_0_198 : _GEN_348; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12355 = 8'hc7 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_350 = ~refillIDX_r & 8'hc7 == req_set ? dirty_0_199 : _GEN_349; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12357 = 8'hc8 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_351 = ~refillIDX_r & 8'hc8 == req_set ? dirty_0_200 : _GEN_350; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12359 = 8'hc9 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_352 = ~refillIDX_r & 8'hc9 == req_set ? dirty_0_201 : _GEN_351; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12361 = 8'hca == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_353 = ~refillIDX_r & 8'hca == req_set ? dirty_0_202 : _GEN_352; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12363 = 8'hcb == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_354 = ~refillIDX_r & 8'hcb == req_set ? dirty_0_203 : _GEN_353; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12365 = 8'hcc == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_355 = ~refillIDX_r & 8'hcc == req_set ? dirty_0_204 : _GEN_354; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12367 = 8'hcd == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_356 = ~refillIDX_r & 8'hcd == req_set ? dirty_0_205 : _GEN_355; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12369 = 8'hce == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_357 = ~refillIDX_r & 8'hce == req_set ? dirty_0_206 : _GEN_356; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12371 = 8'hcf == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_358 = ~refillIDX_r & 8'hcf == req_set ? dirty_0_207 : _GEN_357; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12373 = 8'hd0 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_359 = ~refillIDX_r & 8'hd0 == req_set ? dirty_0_208 : _GEN_358; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12375 = 8'hd1 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_360 = ~refillIDX_r & 8'hd1 == req_set ? dirty_0_209 : _GEN_359; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12377 = 8'hd2 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_361 = ~refillIDX_r & 8'hd2 == req_set ? dirty_0_210 : _GEN_360; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12379 = 8'hd3 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_362 = ~refillIDX_r & 8'hd3 == req_set ? dirty_0_211 : _GEN_361; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12381 = 8'hd4 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_363 = ~refillIDX_r & 8'hd4 == req_set ? dirty_0_212 : _GEN_362; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12383 = 8'hd5 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_364 = ~refillIDX_r & 8'hd5 == req_set ? dirty_0_213 : _GEN_363; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12385 = 8'hd6 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_365 = ~refillIDX_r & 8'hd6 == req_set ? dirty_0_214 : _GEN_364; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12387 = 8'hd7 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_366 = ~refillIDX_r & 8'hd7 == req_set ? dirty_0_215 : _GEN_365; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12389 = 8'hd8 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_367 = ~refillIDX_r & 8'hd8 == req_set ? dirty_0_216 : _GEN_366; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12391 = 8'hd9 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_368 = ~refillIDX_r & 8'hd9 == req_set ? dirty_0_217 : _GEN_367; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12393 = 8'hda == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_369 = ~refillIDX_r & 8'hda == req_set ? dirty_0_218 : _GEN_368; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12395 = 8'hdb == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_370 = ~refillIDX_r & 8'hdb == req_set ? dirty_0_219 : _GEN_369; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12397 = 8'hdc == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_371 = ~refillIDX_r & 8'hdc == req_set ? dirty_0_220 : _GEN_370; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12399 = 8'hdd == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_372 = ~refillIDX_r & 8'hdd == req_set ? dirty_0_221 : _GEN_371; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12401 = 8'hde == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_373 = ~refillIDX_r & 8'hde == req_set ? dirty_0_222 : _GEN_372; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12403 = 8'hdf == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_374 = ~refillIDX_r & 8'hdf == req_set ? dirty_0_223 : _GEN_373; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12405 = 8'he0 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_375 = ~refillIDX_r & 8'he0 == req_set ? dirty_0_224 : _GEN_374; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12407 = 8'he1 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_376 = ~refillIDX_r & 8'he1 == req_set ? dirty_0_225 : _GEN_375; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12409 = 8'he2 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_377 = ~refillIDX_r & 8'he2 == req_set ? dirty_0_226 : _GEN_376; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12411 = 8'he3 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_378 = ~refillIDX_r & 8'he3 == req_set ? dirty_0_227 : _GEN_377; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12413 = 8'he4 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_379 = ~refillIDX_r & 8'he4 == req_set ? dirty_0_228 : _GEN_378; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12415 = 8'he5 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_380 = ~refillIDX_r & 8'he5 == req_set ? dirty_0_229 : _GEN_379; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12417 = 8'he6 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_381 = ~refillIDX_r & 8'he6 == req_set ? dirty_0_230 : _GEN_380; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12419 = 8'he7 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_382 = ~refillIDX_r & 8'he7 == req_set ? dirty_0_231 : _GEN_381; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12421 = 8'he8 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_383 = ~refillIDX_r & 8'he8 == req_set ? dirty_0_232 : _GEN_382; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12423 = 8'he9 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_384 = ~refillIDX_r & 8'he9 == req_set ? dirty_0_233 : _GEN_383; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12425 = 8'hea == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_385 = ~refillIDX_r & 8'hea == req_set ? dirty_0_234 : _GEN_384; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12427 = 8'heb == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_386 = ~refillIDX_r & 8'heb == req_set ? dirty_0_235 : _GEN_385; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12429 = 8'hec == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_387 = ~refillIDX_r & 8'hec == req_set ? dirty_0_236 : _GEN_386; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12431 = 8'hed == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_388 = ~refillIDX_r & 8'hed == req_set ? dirty_0_237 : _GEN_387; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12433 = 8'hee == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_389 = ~refillIDX_r & 8'hee == req_set ? dirty_0_238 : _GEN_388; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12435 = 8'hef == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_390 = ~refillIDX_r & 8'hef == req_set ? dirty_0_239 : _GEN_389; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12437 = 8'hf0 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_391 = ~refillIDX_r & 8'hf0 == req_set ? dirty_0_240 : _GEN_390; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12439 = 8'hf1 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_392 = ~refillIDX_r & 8'hf1 == req_set ? dirty_0_241 : _GEN_391; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12441 = 8'hf2 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_393 = ~refillIDX_r & 8'hf2 == req_set ? dirty_0_242 : _GEN_392; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12443 = 8'hf3 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_394 = ~refillIDX_r & 8'hf3 == req_set ? dirty_0_243 : _GEN_393; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12445 = 8'hf4 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_395 = ~refillIDX_r & 8'hf4 == req_set ? dirty_0_244 : _GEN_394; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12447 = 8'hf5 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_396 = ~refillIDX_r & 8'hf5 == req_set ? dirty_0_245 : _GEN_395; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12449 = 8'hf6 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_397 = ~refillIDX_r & 8'hf6 == req_set ? dirty_0_246 : _GEN_396; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12451 = 8'hf7 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_398 = ~refillIDX_r & 8'hf7 == req_set ? dirty_0_247 : _GEN_397; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12453 = 8'hf8 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_399 = ~refillIDX_r & 8'hf8 == req_set ? dirty_0_248 : _GEN_398; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12455 = 8'hf9 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_400 = ~refillIDX_r & 8'hf9 == req_set ? dirty_0_249 : _GEN_399; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12457 = 8'hfa == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_401 = ~refillIDX_r & 8'hfa == req_set ? dirty_0_250 : _GEN_400; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12459 = 8'hfb == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_402 = ~refillIDX_r & 8'hfb == req_set ? dirty_0_251 : _GEN_401; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12461 = 8'hfc == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_403 = ~refillIDX_r & 8'hfc == req_set ? dirty_0_252 : _GEN_402; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12463 = 8'hfd == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_404 = ~refillIDX_r & 8'hfd == req_set ? dirty_0_253 : _GEN_403; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12465 = 8'hfe == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_405 = ~refillIDX_r & 8'hfe == req_set ? dirty_0_254 : _GEN_404; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12467 = 8'hff == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_406 = ~refillIDX_r & 8'hff == req_set ? dirty_0_255 : _GEN_405; // @[dcache.scala 345:{54,54}]
  wire  _GEN_12468 = 8'h0 == req_set; // @[dcache.scala 345:{54,54}]
  wire  _GEN_407 = refillIDX_r & 8'h0 == req_set ? dirty_1_0 : _GEN_406; // @[dcache.scala 345:{54,54}]
  wire  _GEN_408 = refillIDX_r & 8'h1 == req_set ? dirty_1_1 : _GEN_407; // @[dcache.scala 345:{54,54}]
  wire  _GEN_409 = refillIDX_r & 8'h2 == req_set ? dirty_1_2 : _GEN_408; // @[dcache.scala 345:{54,54}]
  wire  _GEN_410 = refillIDX_r & 8'h3 == req_set ? dirty_1_3 : _GEN_409; // @[dcache.scala 345:{54,54}]
  wire  _GEN_411 = refillIDX_r & 8'h4 == req_set ? dirty_1_4 : _GEN_410; // @[dcache.scala 345:{54,54}]
  wire  _GEN_412 = refillIDX_r & 8'h5 == req_set ? dirty_1_5 : _GEN_411; // @[dcache.scala 345:{54,54}]
  wire  _GEN_413 = refillIDX_r & 8'h6 == req_set ? dirty_1_6 : _GEN_412; // @[dcache.scala 345:{54,54}]
  wire  _GEN_414 = refillIDX_r & 8'h7 == req_set ? dirty_1_7 : _GEN_413; // @[dcache.scala 345:{54,54}]
  wire  _GEN_415 = refillIDX_r & 8'h8 == req_set ? dirty_1_8 : _GEN_414; // @[dcache.scala 345:{54,54}]
  wire  _GEN_416 = refillIDX_r & 8'h9 == req_set ? dirty_1_9 : _GEN_415; // @[dcache.scala 345:{54,54}]
  wire  _GEN_417 = refillIDX_r & 8'ha == req_set ? dirty_1_10 : _GEN_416; // @[dcache.scala 345:{54,54}]
  wire  _GEN_418 = refillIDX_r & 8'hb == req_set ? dirty_1_11 : _GEN_417; // @[dcache.scala 345:{54,54}]
  wire  _GEN_419 = refillIDX_r & 8'hc == req_set ? dirty_1_12 : _GEN_418; // @[dcache.scala 345:{54,54}]
  wire  _GEN_420 = refillIDX_r & 8'hd == req_set ? dirty_1_13 : _GEN_419; // @[dcache.scala 345:{54,54}]
  wire  _GEN_421 = refillIDX_r & 8'he == req_set ? dirty_1_14 : _GEN_420; // @[dcache.scala 345:{54,54}]
  wire  _GEN_422 = refillIDX_r & 8'hf == req_set ? dirty_1_15 : _GEN_421; // @[dcache.scala 345:{54,54}]
  wire  _GEN_423 = refillIDX_r & 8'h10 == req_set ? dirty_1_16 : _GEN_422; // @[dcache.scala 345:{54,54}]
  wire  _GEN_424 = refillIDX_r & 8'h11 == req_set ? dirty_1_17 : _GEN_423; // @[dcache.scala 345:{54,54}]
  wire  _GEN_425 = refillIDX_r & 8'h12 == req_set ? dirty_1_18 : _GEN_424; // @[dcache.scala 345:{54,54}]
  wire  _GEN_426 = refillIDX_r & 8'h13 == req_set ? dirty_1_19 : _GEN_425; // @[dcache.scala 345:{54,54}]
  wire  _GEN_427 = refillIDX_r & 8'h14 == req_set ? dirty_1_20 : _GEN_426; // @[dcache.scala 345:{54,54}]
  wire  _GEN_428 = refillIDX_r & 8'h15 == req_set ? dirty_1_21 : _GEN_427; // @[dcache.scala 345:{54,54}]
  wire  _GEN_429 = refillIDX_r & 8'h16 == req_set ? dirty_1_22 : _GEN_428; // @[dcache.scala 345:{54,54}]
  wire  _GEN_430 = refillIDX_r & 8'h17 == req_set ? dirty_1_23 : _GEN_429; // @[dcache.scala 345:{54,54}]
  wire  _GEN_431 = refillIDX_r & 8'h18 == req_set ? dirty_1_24 : _GEN_430; // @[dcache.scala 345:{54,54}]
  wire  _GEN_432 = refillIDX_r & 8'h19 == req_set ? dirty_1_25 : _GEN_431; // @[dcache.scala 345:{54,54}]
  wire  _GEN_433 = refillIDX_r & 8'h1a == req_set ? dirty_1_26 : _GEN_432; // @[dcache.scala 345:{54,54}]
  wire  _GEN_434 = refillIDX_r & 8'h1b == req_set ? dirty_1_27 : _GEN_433; // @[dcache.scala 345:{54,54}]
  wire  _GEN_435 = refillIDX_r & 8'h1c == req_set ? dirty_1_28 : _GEN_434; // @[dcache.scala 345:{54,54}]
  wire  _GEN_436 = refillIDX_r & 8'h1d == req_set ? dirty_1_29 : _GEN_435; // @[dcache.scala 345:{54,54}]
  wire  _GEN_437 = refillIDX_r & 8'h1e == req_set ? dirty_1_30 : _GEN_436; // @[dcache.scala 345:{54,54}]
  wire  _GEN_438 = refillIDX_r & 8'h1f == req_set ? dirty_1_31 : _GEN_437; // @[dcache.scala 345:{54,54}]
  wire  _GEN_439 = refillIDX_r & 8'h20 == req_set ? dirty_1_32 : _GEN_438; // @[dcache.scala 345:{54,54}]
  wire  _GEN_440 = refillIDX_r & 8'h21 == req_set ? dirty_1_33 : _GEN_439; // @[dcache.scala 345:{54,54}]
  wire  _GEN_441 = refillIDX_r & 8'h22 == req_set ? dirty_1_34 : _GEN_440; // @[dcache.scala 345:{54,54}]
  wire  _GEN_442 = refillIDX_r & 8'h23 == req_set ? dirty_1_35 : _GEN_441; // @[dcache.scala 345:{54,54}]
  wire  _GEN_443 = refillIDX_r & 8'h24 == req_set ? dirty_1_36 : _GEN_442; // @[dcache.scala 345:{54,54}]
  wire  _GEN_444 = refillIDX_r & 8'h25 == req_set ? dirty_1_37 : _GEN_443; // @[dcache.scala 345:{54,54}]
  wire  _GEN_445 = refillIDX_r & 8'h26 == req_set ? dirty_1_38 : _GEN_444; // @[dcache.scala 345:{54,54}]
  wire  _GEN_446 = refillIDX_r & 8'h27 == req_set ? dirty_1_39 : _GEN_445; // @[dcache.scala 345:{54,54}]
  wire  _GEN_447 = refillIDX_r & 8'h28 == req_set ? dirty_1_40 : _GEN_446; // @[dcache.scala 345:{54,54}]
  wire  _GEN_448 = refillIDX_r & 8'h29 == req_set ? dirty_1_41 : _GEN_447; // @[dcache.scala 345:{54,54}]
  wire  _GEN_449 = refillIDX_r & 8'h2a == req_set ? dirty_1_42 : _GEN_448; // @[dcache.scala 345:{54,54}]
  wire  _GEN_450 = refillIDX_r & 8'h2b == req_set ? dirty_1_43 : _GEN_449; // @[dcache.scala 345:{54,54}]
  wire  _GEN_451 = refillIDX_r & 8'h2c == req_set ? dirty_1_44 : _GEN_450; // @[dcache.scala 345:{54,54}]
  wire  _GEN_452 = refillIDX_r & 8'h2d == req_set ? dirty_1_45 : _GEN_451; // @[dcache.scala 345:{54,54}]
  wire  _GEN_453 = refillIDX_r & 8'h2e == req_set ? dirty_1_46 : _GEN_452; // @[dcache.scala 345:{54,54}]
  wire  _GEN_454 = refillIDX_r & 8'h2f == req_set ? dirty_1_47 : _GEN_453; // @[dcache.scala 345:{54,54}]
  wire  _GEN_455 = refillIDX_r & 8'h30 == req_set ? dirty_1_48 : _GEN_454; // @[dcache.scala 345:{54,54}]
  wire  _GEN_456 = refillIDX_r & 8'h31 == req_set ? dirty_1_49 : _GEN_455; // @[dcache.scala 345:{54,54}]
  wire  _GEN_457 = refillIDX_r & 8'h32 == req_set ? dirty_1_50 : _GEN_456; // @[dcache.scala 345:{54,54}]
  wire  _GEN_458 = refillIDX_r & 8'h33 == req_set ? dirty_1_51 : _GEN_457; // @[dcache.scala 345:{54,54}]
  wire  _GEN_459 = refillIDX_r & 8'h34 == req_set ? dirty_1_52 : _GEN_458; // @[dcache.scala 345:{54,54}]
  wire  _GEN_460 = refillIDX_r & 8'h35 == req_set ? dirty_1_53 : _GEN_459; // @[dcache.scala 345:{54,54}]
  wire  _GEN_461 = refillIDX_r & 8'h36 == req_set ? dirty_1_54 : _GEN_460; // @[dcache.scala 345:{54,54}]
  wire  _GEN_462 = refillIDX_r & 8'h37 == req_set ? dirty_1_55 : _GEN_461; // @[dcache.scala 345:{54,54}]
  wire  _GEN_463 = refillIDX_r & 8'h38 == req_set ? dirty_1_56 : _GEN_462; // @[dcache.scala 345:{54,54}]
  wire  _GEN_464 = refillIDX_r & 8'h39 == req_set ? dirty_1_57 : _GEN_463; // @[dcache.scala 345:{54,54}]
  wire  _GEN_465 = refillIDX_r & 8'h3a == req_set ? dirty_1_58 : _GEN_464; // @[dcache.scala 345:{54,54}]
  wire  _GEN_466 = refillIDX_r & 8'h3b == req_set ? dirty_1_59 : _GEN_465; // @[dcache.scala 345:{54,54}]
  wire  _GEN_467 = refillIDX_r & 8'h3c == req_set ? dirty_1_60 : _GEN_466; // @[dcache.scala 345:{54,54}]
  wire  _GEN_468 = refillIDX_r & 8'h3d == req_set ? dirty_1_61 : _GEN_467; // @[dcache.scala 345:{54,54}]
  wire  _GEN_469 = refillIDX_r & 8'h3e == req_set ? dirty_1_62 : _GEN_468; // @[dcache.scala 345:{54,54}]
  wire  _GEN_470 = refillIDX_r & 8'h3f == req_set ? dirty_1_63 : _GEN_469; // @[dcache.scala 345:{54,54}]
  wire  _GEN_471 = refillIDX_r & 8'h40 == req_set ? dirty_1_64 : _GEN_470; // @[dcache.scala 345:{54,54}]
  wire  _GEN_472 = refillIDX_r & 8'h41 == req_set ? dirty_1_65 : _GEN_471; // @[dcache.scala 345:{54,54}]
  wire  _GEN_473 = refillIDX_r & 8'h42 == req_set ? dirty_1_66 : _GEN_472; // @[dcache.scala 345:{54,54}]
  wire  _GEN_474 = refillIDX_r & 8'h43 == req_set ? dirty_1_67 : _GEN_473; // @[dcache.scala 345:{54,54}]
  wire  _GEN_475 = refillIDX_r & 8'h44 == req_set ? dirty_1_68 : _GEN_474; // @[dcache.scala 345:{54,54}]
  wire  _GEN_476 = refillIDX_r & 8'h45 == req_set ? dirty_1_69 : _GEN_475; // @[dcache.scala 345:{54,54}]
  wire  _GEN_477 = refillIDX_r & 8'h46 == req_set ? dirty_1_70 : _GEN_476; // @[dcache.scala 345:{54,54}]
  wire  _GEN_478 = refillIDX_r & 8'h47 == req_set ? dirty_1_71 : _GEN_477; // @[dcache.scala 345:{54,54}]
  wire  _GEN_479 = refillIDX_r & 8'h48 == req_set ? dirty_1_72 : _GEN_478; // @[dcache.scala 345:{54,54}]
  wire  _GEN_480 = refillIDX_r & 8'h49 == req_set ? dirty_1_73 : _GEN_479; // @[dcache.scala 345:{54,54}]
  wire  _GEN_481 = refillIDX_r & 8'h4a == req_set ? dirty_1_74 : _GEN_480; // @[dcache.scala 345:{54,54}]
  wire  _GEN_482 = refillIDX_r & 8'h4b == req_set ? dirty_1_75 : _GEN_481; // @[dcache.scala 345:{54,54}]
  wire  _GEN_483 = refillIDX_r & 8'h4c == req_set ? dirty_1_76 : _GEN_482; // @[dcache.scala 345:{54,54}]
  wire  _GEN_484 = refillIDX_r & 8'h4d == req_set ? dirty_1_77 : _GEN_483; // @[dcache.scala 345:{54,54}]
  wire  _GEN_485 = refillIDX_r & 8'h4e == req_set ? dirty_1_78 : _GEN_484; // @[dcache.scala 345:{54,54}]
  wire  _GEN_486 = refillIDX_r & 8'h4f == req_set ? dirty_1_79 : _GEN_485; // @[dcache.scala 345:{54,54}]
  wire  _GEN_487 = refillIDX_r & 8'h50 == req_set ? dirty_1_80 : _GEN_486; // @[dcache.scala 345:{54,54}]
  wire  _GEN_488 = refillIDX_r & 8'h51 == req_set ? dirty_1_81 : _GEN_487; // @[dcache.scala 345:{54,54}]
  wire  _GEN_489 = refillIDX_r & 8'h52 == req_set ? dirty_1_82 : _GEN_488; // @[dcache.scala 345:{54,54}]
  wire  _GEN_490 = refillIDX_r & 8'h53 == req_set ? dirty_1_83 : _GEN_489; // @[dcache.scala 345:{54,54}]
  wire  _GEN_491 = refillIDX_r & 8'h54 == req_set ? dirty_1_84 : _GEN_490; // @[dcache.scala 345:{54,54}]
  wire  _GEN_492 = refillIDX_r & 8'h55 == req_set ? dirty_1_85 : _GEN_491; // @[dcache.scala 345:{54,54}]
  wire  _GEN_493 = refillIDX_r & 8'h56 == req_set ? dirty_1_86 : _GEN_492; // @[dcache.scala 345:{54,54}]
  wire  _GEN_494 = refillIDX_r & 8'h57 == req_set ? dirty_1_87 : _GEN_493; // @[dcache.scala 345:{54,54}]
  wire  _GEN_495 = refillIDX_r & 8'h58 == req_set ? dirty_1_88 : _GEN_494; // @[dcache.scala 345:{54,54}]
  wire  _GEN_496 = refillIDX_r & 8'h59 == req_set ? dirty_1_89 : _GEN_495; // @[dcache.scala 345:{54,54}]
  wire  _GEN_497 = refillIDX_r & 8'h5a == req_set ? dirty_1_90 : _GEN_496; // @[dcache.scala 345:{54,54}]
  wire  _GEN_498 = refillIDX_r & 8'h5b == req_set ? dirty_1_91 : _GEN_497; // @[dcache.scala 345:{54,54}]
  wire  _GEN_499 = refillIDX_r & 8'h5c == req_set ? dirty_1_92 : _GEN_498; // @[dcache.scala 345:{54,54}]
  wire  _GEN_500 = refillIDX_r & 8'h5d == req_set ? dirty_1_93 : _GEN_499; // @[dcache.scala 345:{54,54}]
  wire  _GEN_501 = refillIDX_r & 8'h5e == req_set ? dirty_1_94 : _GEN_500; // @[dcache.scala 345:{54,54}]
  wire  _GEN_502 = refillIDX_r & 8'h5f == req_set ? dirty_1_95 : _GEN_501; // @[dcache.scala 345:{54,54}]
  wire  _GEN_503 = refillIDX_r & 8'h60 == req_set ? dirty_1_96 : _GEN_502; // @[dcache.scala 345:{54,54}]
  wire  _GEN_504 = refillIDX_r & 8'h61 == req_set ? dirty_1_97 : _GEN_503; // @[dcache.scala 345:{54,54}]
  wire  _GEN_505 = refillIDX_r & 8'h62 == req_set ? dirty_1_98 : _GEN_504; // @[dcache.scala 345:{54,54}]
  wire  _GEN_506 = refillIDX_r & 8'h63 == req_set ? dirty_1_99 : _GEN_505; // @[dcache.scala 345:{54,54}]
  wire  _GEN_507 = refillIDX_r & 8'h64 == req_set ? dirty_1_100 : _GEN_506; // @[dcache.scala 345:{54,54}]
  wire  _GEN_508 = refillIDX_r & 8'h65 == req_set ? dirty_1_101 : _GEN_507; // @[dcache.scala 345:{54,54}]
  wire  _GEN_509 = refillIDX_r & 8'h66 == req_set ? dirty_1_102 : _GEN_508; // @[dcache.scala 345:{54,54}]
  wire  _GEN_510 = refillIDX_r & 8'h67 == req_set ? dirty_1_103 : _GEN_509; // @[dcache.scala 345:{54,54}]
  wire  _GEN_511 = refillIDX_r & 8'h68 == req_set ? dirty_1_104 : _GEN_510; // @[dcache.scala 345:{54,54}]
  wire  _GEN_512 = refillIDX_r & 8'h69 == req_set ? dirty_1_105 : _GEN_511; // @[dcache.scala 345:{54,54}]
  wire  _GEN_513 = refillIDX_r & 8'h6a == req_set ? dirty_1_106 : _GEN_512; // @[dcache.scala 345:{54,54}]
  wire  _GEN_514 = refillIDX_r & 8'h6b == req_set ? dirty_1_107 : _GEN_513; // @[dcache.scala 345:{54,54}]
  wire  _GEN_515 = refillIDX_r & 8'h6c == req_set ? dirty_1_108 : _GEN_514; // @[dcache.scala 345:{54,54}]
  wire  _GEN_516 = refillIDX_r & 8'h6d == req_set ? dirty_1_109 : _GEN_515; // @[dcache.scala 345:{54,54}]
  wire  _GEN_517 = refillIDX_r & 8'h6e == req_set ? dirty_1_110 : _GEN_516; // @[dcache.scala 345:{54,54}]
  wire  _GEN_518 = refillIDX_r & 8'h6f == req_set ? dirty_1_111 : _GEN_517; // @[dcache.scala 345:{54,54}]
  wire  _GEN_519 = refillIDX_r & 8'h70 == req_set ? dirty_1_112 : _GEN_518; // @[dcache.scala 345:{54,54}]
  wire  _GEN_520 = refillIDX_r & 8'h71 == req_set ? dirty_1_113 : _GEN_519; // @[dcache.scala 345:{54,54}]
  wire  _GEN_521 = refillIDX_r & 8'h72 == req_set ? dirty_1_114 : _GEN_520; // @[dcache.scala 345:{54,54}]
  wire  _GEN_522 = refillIDX_r & 8'h73 == req_set ? dirty_1_115 : _GEN_521; // @[dcache.scala 345:{54,54}]
  wire  _GEN_523 = refillIDX_r & 8'h74 == req_set ? dirty_1_116 : _GEN_522; // @[dcache.scala 345:{54,54}]
  wire  _GEN_524 = refillIDX_r & 8'h75 == req_set ? dirty_1_117 : _GEN_523; // @[dcache.scala 345:{54,54}]
  wire  _GEN_525 = refillIDX_r & 8'h76 == req_set ? dirty_1_118 : _GEN_524; // @[dcache.scala 345:{54,54}]
  wire  _GEN_526 = refillIDX_r & 8'h77 == req_set ? dirty_1_119 : _GEN_525; // @[dcache.scala 345:{54,54}]
  wire  _GEN_527 = refillIDX_r & 8'h78 == req_set ? dirty_1_120 : _GEN_526; // @[dcache.scala 345:{54,54}]
  wire  _GEN_528 = refillIDX_r & 8'h79 == req_set ? dirty_1_121 : _GEN_527; // @[dcache.scala 345:{54,54}]
  wire  _GEN_529 = refillIDX_r & 8'h7a == req_set ? dirty_1_122 : _GEN_528; // @[dcache.scala 345:{54,54}]
  wire  _GEN_530 = refillIDX_r & 8'h7b == req_set ? dirty_1_123 : _GEN_529; // @[dcache.scala 345:{54,54}]
  wire  _GEN_531 = refillIDX_r & 8'h7c == req_set ? dirty_1_124 : _GEN_530; // @[dcache.scala 345:{54,54}]
  wire  _GEN_532 = refillIDX_r & 8'h7d == req_set ? dirty_1_125 : _GEN_531; // @[dcache.scala 345:{54,54}]
  wire  _GEN_533 = refillIDX_r & 8'h7e == req_set ? dirty_1_126 : _GEN_532; // @[dcache.scala 345:{54,54}]
  wire  _GEN_534 = refillIDX_r & 8'h7f == req_set ? dirty_1_127 : _GEN_533; // @[dcache.scala 345:{54,54}]
  wire  _GEN_535 = refillIDX_r & 8'h80 == req_set ? dirty_1_128 : _GEN_534; // @[dcache.scala 345:{54,54}]
  wire  _GEN_536 = refillIDX_r & 8'h81 == req_set ? dirty_1_129 : _GEN_535; // @[dcache.scala 345:{54,54}]
  wire  _GEN_537 = refillIDX_r & 8'h82 == req_set ? dirty_1_130 : _GEN_536; // @[dcache.scala 345:{54,54}]
  wire  _GEN_538 = refillIDX_r & 8'h83 == req_set ? dirty_1_131 : _GEN_537; // @[dcache.scala 345:{54,54}]
  wire  _GEN_539 = refillIDX_r & 8'h84 == req_set ? dirty_1_132 : _GEN_538; // @[dcache.scala 345:{54,54}]
  wire  _GEN_540 = refillIDX_r & 8'h85 == req_set ? dirty_1_133 : _GEN_539; // @[dcache.scala 345:{54,54}]
  wire  _GEN_541 = refillIDX_r & 8'h86 == req_set ? dirty_1_134 : _GEN_540; // @[dcache.scala 345:{54,54}]
  wire  _GEN_542 = refillIDX_r & 8'h87 == req_set ? dirty_1_135 : _GEN_541; // @[dcache.scala 345:{54,54}]
  wire  _GEN_543 = refillIDX_r & 8'h88 == req_set ? dirty_1_136 : _GEN_542; // @[dcache.scala 345:{54,54}]
  wire  _GEN_544 = refillIDX_r & 8'h89 == req_set ? dirty_1_137 : _GEN_543; // @[dcache.scala 345:{54,54}]
  wire  _GEN_545 = refillIDX_r & 8'h8a == req_set ? dirty_1_138 : _GEN_544; // @[dcache.scala 345:{54,54}]
  wire  _GEN_546 = refillIDX_r & 8'h8b == req_set ? dirty_1_139 : _GEN_545; // @[dcache.scala 345:{54,54}]
  wire  _GEN_547 = refillIDX_r & 8'h8c == req_set ? dirty_1_140 : _GEN_546; // @[dcache.scala 345:{54,54}]
  wire  _GEN_548 = refillIDX_r & 8'h8d == req_set ? dirty_1_141 : _GEN_547; // @[dcache.scala 345:{54,54}]
  wire  _GEN_549 = refillIDX_r & 8'h8e == req_set ? dirty_1_142 : _GEN_548; // @[dcache.scala 345:{54,54}]
  wire  _GEN_550 = refillIDX_r & 8'h8f == req_set ? dirty_1_143 : _GEN_549; // @[dcache.scala 345:{54,54}]
  wire  _GEN_551 = refillIDX_r & 8'h90 == req_set ? dirty_1_144 : _GEN_550; // @[dcache.scala 345:{54,54}]
  wire  _GEN_552 = refillIDX_r & 8'h91 == req_set ? dirty_1_145 : _GEN_551; // @[dcache.scala 345:{54,54}]
  wire  _GEN_553 = refillIDX_r & 8'h92 == req_set ? dirty_1_146 : _GEN_552; // @[dcache.scala 345:{54,54}]
  wire  _GEN_554 = refillIDX_r & 8'h93 == req_set ? dirty_1_147 : _GEN_553; // @[dcache.scala 345:{54,54}]
  wire  _GEN_555 = refillIDX_r & 8'h94 == req_set ? dirty_1_148 : _GEN_554; // @[dcache.scala 345:{54,54}]
  wire  _GEN_556 = refillIDX_r & 8'h95 == req_set ? dirty_1_149 : _GEN_555; // @[dcache.scala 345:{54,54}]
  wire  _GEN_557 = refillIDX_r & 8'h96 == req_set ? dirty_1_150 : _GEN_556; // @[dcache.scala 345:{54,54}]
  wire  _GEN_558 = refillIDX_r & 8'h97 == req_set ? dirty_1_151 : _GEN_557; // @[dcache.scala 345:{54,54}]
  wire  _GEN_559 = refillIDX_r & 8'h98 == req_set ? dirty_1_152 : _GEN_558; // @[dcache.scala 345:{54,54}]
  wire  _GEN_560 = refillIDX_r & 8'h99 == req_set ? dirty_1_153 : _GEN_559; // @[dcache.scala 345:{54,54}]
  wire  _GEN_561 = refillIDX_r & 8'h9a == req_set ? dirty_1_154 : _GEN_560; // @[dcache.scala 345:{54,54}]
  wire  _GEN_562 = refillIDX_r & 8'h9b == req_set ? dirty_1_155 : _GEN_561; // @[dcache.scala 345:{54,54}]
  wire  _GEN_563 = refillIDX_r & 8'h9c == req_set ? dirty_1_156 : _GEN_562; // @[dcache.scala 345:{54,54}]
  wire  _GEN_564 = refillIDX_r & 8'h9d == req_set ? dirty_1_157 : _GEN_563; // @[dcache.scala 345:{54,54}]
  wire  _GEN_565 = refillIDX_r & 8'h9e == req_set ? dirty_1_158 : _GEN_564; // @[dcache.scala 345:{54,54}]
  wire  _GEN_566 = refillIDX_r & 8'h9f == req_set ? dirty_1_159 : _GEN_565; // @[dcache.scala 345:{54,54}]
  wire  _GEN_567 = refillIDX_r & 8'ha0 == req_set ? dirty_1_160 : _GEN_566; // @[dcache.scala 345:{54,54}]
  wire  _GEN_568 = refillIDX_r & 8'ha1 == req_set ? dirty_1_161 : _GEN_567; // @[dcache.scala 345:{54,54}]
  wire  _GEN_569 = refillIDX_r & 8'ha2 == req_set ? dirty_1_162 : _GEN_568; // @[dcache.scala 345:{54,54}]
  wire  _GEN_570 = refillIDX_r & 8'ha3 == req_set ? dirty_1_163 : _GEN_569; // @[dcache.scala 345:{54,54}]
  wire  _GEN_571 = refillIDX_r & 8'ha4 == req_set ? dirty_1_164 : _GEN_570; // @[dcache.scala 345:{54,54}]
  wire  _GEN_572 = refillIDX_r & 8'ha5 == req_set ? dirty_1_165 : _GEN_571; // @[dcache.scala 345:{54,54}]
  wire  _GEN_573 = refillIDX_r & 8'ha6 == req_set ? dirty_1_166 : _GEN_572; // @[dcache.scala 345:{54,54}]
  wire  _GEN_574 = refillIDX_r & 8'ha7 == req_set ? dirty_1_167 : _GEN_573; // @[dcache.scala 345:{54,54}]
  wire  _GEN_575 = refillIDX_r & 8'ha8 == req_set ? dirty_1_168 : _GEN_574; // @[dcache.scala 345:{54,54}]
  wire  _GEN_576 = refillIDX_r & 8'ha9 == req_set ? dirty_1_169 : _GEN_575; // @[dcache.scala 345:{54,54}]
  wire  _GEN_577 = refillIDX_r & 8'haa == req_set ? dirty_1_170 : _GEN_576; // @[dcache.scala 345:{54,54}]
  wire  _GEN_578 = refillIDX_r & 8'hab == req_set ? dirty_1_171 : _GEN_577; // @[dcache.scala 345:{54,54}]
  wire  _GEN_579 = refillIDX_r & 8'hac == req_set ? dirty_1_172 : _GEN_578; // @[dcache.scala 345:{54,54}]
  wire  _GEN_580 = refillIDX_r & 8'had == req_set ? dirty_1_173 : _GEN_579; // @[dcache.scala 345:{54,54}]
  wire  _GEN_581 = refillIDX_r & 8'hae == req_set ? dirty_1_174 : _GEN_580; // @[dcache.scala 345:{54,54}]
  wire  _GEN_582 = refillIDX_r & 8'haf == req_set ? dirty_1_175 : _GEN_581; // @[dcache.scala 345:{54,54}]
  wire  _GEN_583 = refillIDX_r & 8'hb0 == req_set ? dirty_1_176 : _GEN_582; // @[dcache.scala 345:{54,54}]
  wire  _GEN_584 = refillIDX_r & 8'hb1 == req_set ? dirty_1_177 : _GEN_583; // @[dcache.scala 345:{54,54}]
  wire  _GEN_585 = refillIDX_r & 8'hb2 == req_set ? dirty_1_178 : _GEN_584; // @[dcache.scala 345:{54,54}]
  wire  _GEN_586 = refillIDX_r & 8'hb3 == req_set ? dirty_1_179 : _GEN_585; // @[dcache.scala 345:{54,54}]
  wire  _GEN_587 = refillIDX_r & 8'hb4 == req_set ? dirty_1_180 : _GEN_586; // @[dcache.scala 345:{54,54}]
  wire  _GEN_588 = refillIDX_r & 8'hb5 == req_set ? dirty_1_181 : _GEN_587; // @[dcache.scala 345:{54,54}]
  wire  _GEN_589 = refillIDX_r & 8'hb6 == req_set ? dirty_1_182 : _GEN_588; // @[dcache.scala 345:{54,54}]
  wire  _GEN_590 = refillIDX_r & 8'hb7 == req_set ? dirty_1_183 : _GEN_589; // @[dcache.scala 345:{54,54}]
  wire  _GEN_591 = refillIDX_r & 8'hb8 == req_set ? dirty_1_184 : _GEN_590; // @[dcache.scala 345:{54,54}]
  wire  _GEN_592 = refillIDX_r & 8'hb9 == req_set ? dirty_1_185 : _GEN_591; // @[dcache.scala 345:{54,54}]
  wire  _GEN_593 = refillIDX_r & 8'hba == req_set ? dirty_1_186 : _GEN_592; // @[dcache.scala 345:{54,54}]
  wire  _GEN_594 = refillIDX_r & 8'hbb == req_set ? dirty_1_187 : _GEN_593; // @[dcache.scala 345:{54,54}]
  wire  _GEN_595 = refillIDX_r & 8'hbc == req_set ? dirty_1_188 : _GEN_594; // @[dcache.scala 345:{54,54}]
  wire  _GEN_596 = refillIDX_r & 8'hbd == req_set ? dirty_1_189 : _GEN_595; // @[dcache.scala 345:{54,54}]
  wire  _GEN_597 = refillIDX_r & 8'hbe == req_set ? dirty_1_190 : _GEN_596; // @[dcache.scala 345:{54,54}]
  wire  _GEN_598 = refillIDX_r & 8'hbf == req_set ? dirty_1_191 : _GEN_597; // @[dcache.scala 345:{54,54}]
  wire  _GEN_599 = refillIDX_r & 8'hc0 == req_set ? dirty_1_192 : _GEN_598; // @[dcache.scala 345:{54,54}]
  wire  _GEN_600 = refillIDX_r & 8'hc1 == req_set ? dirty_1_193 : _GEN_599; // @[dcache.scala 345:{54,54}]
  wire  _GEN_601 = refillIDX_r & 8'hc2 == req_set ? dirty_1_194 : _GEN_600; // @[dcache.scala 345:{54,54}]
  wire  _GEN_602 = refillIDX_r & 8'hc3 == req_set ? dirty_1_195 : _GEN_601; // @[dcache.scala 345:{54,54}]
  wire  _GEN_603 = refillIDX_r & 8'hc4 == req_set ? dirty_1_196 : _GEN_602; // @[dcache.scala 345:{54,54}]
  wire  _GEN_604 = refillIDX_r & 8'hc5 == req_set ? dirty_1_197 : _GEN_603; // @[dcache.scala 345:{54,54}]
  wire  _GEN_605 = refillIDX_r & 8'hc6 == req_set ? dirty_1_198 : _GEN_604; // @[dcache.scala 345:{54,54}]
  wire  _GEN_606 = refillIDX_r & 8'hc7 == req_set ? dirty_1_199 : _GEN_605; // @[dcache.scala 345:{54,54}]
  wire  _GEN_607 = refillIDX_r & 8'hc8 == req_set ? dirty_1_200 : _GEN_606; // @[dcache.scala 345:{54,54}]
  wire  _GEN_608 = refillIDX_r & 8'hc9 == req_set ? dirty_1_201 : _GEN_607; // @[dcache.scala 345:{54,54}]
  wire  _GEN_609 = refillIDX_r & 8'hca == req_set ? dirty_1_202 : _GEN_608; // @[dcache.scala 345:{54,54}]
  wire  _GEN_610 = refillIDX_r & 8'hcb == req_set ? dirty_1_203 : _GEN_609; // @[dcache.scala 345:{54,54}]
  wire  _GEN_611 = refillIDX_r & 8'hcc == req_set ? dirty_1_204 : _GEN_610; // @[dcache.scala 345:{54,54}]
  wire  _GEN_612 = refillIDX_r & 8'hcd == req_set ? dirty_1_205 : _GEN_611; // @[dcache.scala 345:{54,54}]
  wire  _GEN_613 = refillIDX_r & 8'hce == req_set ? dirty_1_206 : _GEN_612; // @[dcache.scala 345:{54,54}]
  wire  _GEN_614 = refillIDX_r & 8'hcf == req_set ? dirty_1_207 : _GEN_613; // @[dcache.scala 345:{54,54}]
  wire  _GEN_615 = refillIDX_r & 8'hd0 == req_set ? dirty_1_208 : _GEN_614; // @[dcache.scala 345:{54,54}]
  wire  _GEN_616 = refillIDX_r & 8'hd1 == req_set ? dirty_1_209 : _GEN_615; // @[dcache.scala 345:{54,54}]
  wire  _GEN_617 = refillIDX_r & 8'hd2 == req_set ? dirty_1_210 : _GEN_616; // @[dcache.scala 345:{54,54}]
  wire  _GEN_618 = refillIDX_r & 8'hd3 == req_set ? dirty_1_211 : _GEN_617; // @[dcache.scala 345:{54,54}]
  wire  _GEN_619 = refillIDX_r & 8'hd4 == req_set ? dirty_1_212 : _GEN_618; // @[dcache.scala 345:{54,54}]
  wire  _GEN_620 = refillIDX_r & 8'hd5 == req_set ? dirty_1_213 : _GEN_619; // @[dcache.scala 345:{54,54}]
  wire  _GEN_621 = refillIDX_r & 8'hd6 == req_set ? dirty_1_214 : _GEN_620; // @[dcache.scala 345:{54,54}]
  wire  _GEN_622 = refillIDX_r & 8'hd7 == req_set ? dirty_1_215 : _GEN_621; // @[dcache.scala 345:{54,54}]
  wire  _GEN_623 = refillIDX_r & 8'hd8 == req_set ? dirty_1_216 : _GEN_622; // @[dcache.scala 345:{54,54}]
  wire  _GEN_624 = refillIDX_r & 8'hd9 == req_set ? dirty_1_217 : _GEN_623; // @[dcache.scala 345:{54,54}]
  wire  _GEN_625 = refillIDX_r & 8'hda == req_set ? dirty_1_218 : _GEN_624; // @[dcache.scala 345:{54,54}]
  wire  _GEN_626 = refillIDX_r & 8'hdb == req_set ? dirty_1_219 : _GEN_625; // @[dcache.scala 345:{54,54}]
  wire  _GEN_627 = refillIDX_r & 8'hdc == req_set ? dirty_1_220 : _GEN_626; // @[dcache.scala 345:{54,54}]
  wire  _GEN_628 = refillIDX_r & 8'hdd == req_set ? dirty_1_221 : _GEN_627; // @[dcache.scala 345:{54,54}]
  wire  _GEN_629 = refillIDX_r & 8'hde == req_set ? dirty_1_222 : _GEN_628; // @[dcache.scala 345:{54,54}]
  wire  _GEN_630 = refillIDX_r & 8'hdf == req_set ? dirty_1_223 : _GEN_629; // @[dcache.scala 345:{54,54}]
  wire  _GEN_631 = refillIDX_r & 8'he0 == req_set ? dirty_1_224 : _GEN_630; // @[dcache.scala 345:{54,54}]
  wire  _GEN_632 = refillIDX_r & 8'he1 == req_set ? dirty_1_225 : _GEN_631; // @[dcache.scala 345:{54,54}]
  wire  _GEN_633 = refillIDX_r & 8'he2 == req_set ? dirty_1_226 : _GEN_632; // @[dcache.scala 345:{54,54}]
  wire  _GEN_634 = refillIDX_r & 8'he3 == req_set ? dirty_1_227 : _GEN_633; // @[dcache.scala 345:{54,54}]
  wire  _GEN_635 = refillIDX_r & 8'he4 == req_set ? dirty_1_228 : _GEN_634; // @[dcache.scala 345:{54,54}]
  wire  _GEN_636 = refillIDX_r & 8'he5 == req_set ? dirty_1_229 : _GEN_635; // @[dcache.scala 345:{54,54}]
  wire  _GEN_637 = refillIDX_r & 8'he6 == req_set ? dirty_1_230 : _GEN_636; // @[dcache.scala 345:{54,54}]
  wire  _GEN_638 = refillIDX_r & 8'he7 == req_set ? dirty_1_231 : _GEN_637; // @[dcache.scala 345:{54,54}]
  wire  _GEN_639 = refillIDX_r & 8'he8 == req_set ? dirty_1_232 : _GEN_638; // @[dcache.scala 345:{54,54}]
  wire  _GEN_640 = refillIDX_r & 8'he9 == req_set ? dirty_1_233 : _GEN_639; // @[dcache.scala 345:{54,54}]
  wire  _GEN_641 = refillIDX_r & 8'hea == req_set ? dirty_1_234 : _GEN_640; // @[dcache.scala 345:{54,54}]
  wire  _GEN_642 = refillIDX_r & 8'heb == req_set ? dirty_1_235 : _GEN_641; // @[dcache.scala 345:{54,54}]
  wire  _GEN_643 = refillIDX_r & 8'hec == req_set ? dirty_1_236 : _GEN_642; // @[dcache.scala 345:{54,54}]
  wire  _GEN_644 = refillIDX_r & 8'hed == req_set ? dirty_1_237 : _GEN_643; // @[dcache.scala 345:{54,54}]
  wire  _GEN_645 = refillIDX_r & 8'hee == req_set ? dirty_1_238 : _GEN_644; // @[dcache.scala 345:{54,54}]
  wire  _GEN_646 = refillIDX_r & 8'hef == req_set ? dirty_1_239 : _GEN_645; // @[dcache.scala 345:{54,54}]
  wire  _GEN_647 = refillIDX_r & 8'hf0 == req_set ? dirty_1_240 : _GEN_646; // @[dcache.scala 345:{54,54}]
  wire  _GEN_648 = refillIDX_r & 8'hf1 == req_set ? dirty_1_241 : _GEN_647; // @[dcache.scala 345:{54,54}]
  wire  _GEN_649 = refillIDX_r & 8'hf2 == req_set ? dirty_1_242 : _GEN_648; // @[dcache.scala 345:{54,54}]
  wire  _GEN_650 = refillIDX_r & 8'hf3 == req_set ? dirty_1_243 : _GEN_649; // @[dcache.scala 345:{54,54}]
  wire  _GEN_651 = refillIDX_r & 8'hf4 == req_set ? dirty_1_244 : _GEN_650; // @[dcache.scala 345:{54,54}]
  wire  _GEN_652 = refillIDX_r & 8'hf5 == req_set ? dirty_1_245 : _GEN_651; // @[dcache.scala 345:{54,54}]
  wire  _GEN_653 = refillIDX_r & 8'hf6 == req_set ? dirty_1_246 : _GEN_652; // @[dcache.scala 345:{54,54}]
  wire  _GEN_654 = refillIDX_r & 8'hf7 == req_set ? dirty_1_247 : _GEN_653; // @[dcache.scala 345:{54,54}]
  wire  _GEN_655 = refillIDX_r & 8'hf8 == req_set ? dirty_1_248 : _GEN_654; // @[dcache.scala 345:{54,54}]
  wire  _GEN_656 = refillIDX_r & 8'hf9 == req_set ? dirty_1_249 : _GEN_655; // @[dcache.scala 345:{54,54}]
  wire  _GEN_657 = refillIDX_r & 8'hfa == req_set ? dirty_1_250 : _GEN_656; // @[dcache.scala 345:{54,54}]
  wire  _GEN_658 = refillIDX_r & 8'hfb == req_set ? dirty_1_251 : _GEN_657; // @[dcache.scala 345:{54,54}]
  wire  _GEN_659 = refillIDX_r & 8'hfc == req_set ? dirty_1_252 : _GEN_658; // @[dcache.scala 345:{54,54}]
  wire  _GEN_660 = refillIDX_r & 8'hfd == req_set ? dirty_1_253 : _GEN_659; // @[dcache.scala 345:{54,54}]
  wire  _GEN_661 = refillIDX_r & 8'hfe == req_set ? dirty_1_254 : _GEN_660; // @[dcache.scala 345:{54,54}]
  wire  _GEN_662 = refillIDX_r & 8'hff == req_set ? dirty_1_255 : _GEN_661; // @[dcache.scala 345:{54,54}]
  wire [20:0] _GEN_664 = refillIDX_r ? tagv_r_1 : tagv_r_0; // @[dcache.scala 347:{67,67}]
  wire [31:0] _wr_addr_T_1 = {_GEN_664[19:0],req_set,4'h0}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_666 = refillIDX_r ? data_1_1_douta : data_0_1_douta; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_668 = refillIDX_r ? data_1_0_douta : data_0_0_douta; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_670 = refillIDX_r ? data_1_3_douta : data_0_3_douta; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_672 = refillIDX_r ? data_1_2_douta : data_0_2_douta; // @[Cat.scala 33:{92,92}]
  wire [127:0] _wr_data_T = {_GEN_670,_GEN_672,_GEN_666,_GEN_668}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_674 = _GEN_662 ? _wr_addr_T_1 : 32'h0; // @[dcache.scala 163:25 345:54 347:37]
  wire [127:0] _GEN_675 = _GEN_662 ? _wr_data_T : 128'h0; // @[dcache.scala 165:25 345:54 348:37]
  wire [2:0] _GEN_676 = _GEN_662 ? 3'h4 : 3'h0; // @[dcache.scala 162:25 345:54 350:37]
  wire [3:0] _GEN_677 = _GEN_662 ? 4'hf : 4'h0; // @[dcache.scala 164:25 345:54 351:37]
  wire  _T_43 = req_op & req_uncached; // @[dcache.scala 354:34]
  wire [31:0] _wr_addr_T_2 = {req_tag,req_set,req_offset}; // @[Cat.scala 33:92]
  wire [127:0] _wr_data_T_1 = {96'h0,req_wdata_0}; // @[Cat.scala 33:92]
  wire [2:0] _wr_type_T = {{1'd0}, req_lstype[2:1]}; // @[dcache.scala 360:47]
  wire [2:0] _GEN_678 = req_op & req_uncached ? 3'h0 : 3'h3; // @[dcache.scala 334:23 354:51 355:33]
  wire [31:0] _GEN_680 = req_op & req_uncached ? _wr_addr_T_2 : 32'h0; // @[dcache.scala 163:25 354:51 357:33]
  wire [127:0] _GEN_681 = req_op & req_uncached ? _wr_data_T_1 : 128'h0; // @[dcache.scala 165:25 354:51 358:33]
  wire [3:0] _GEN_682 = req_op & req_uncached ? req_wstrb_0 : 4'h0; // @[dcache.scala 164:25 354:51 359:33]
  wire [2:0] _GEN_683 = req_op & req_uncached ? _wr_type_T : 3'h0; // @[dcache.scala 162:25 354:51 360:33]
  wire [2:0] _GEN_684 = _hit_T | writeBack ? 3'h4 : _GEN_678; // @[dcache.scala 343:55 344:37]
  wire  _GEN_685 = _hit_T | writeBack ? _GEN_662 : _T_43; // @[dcache.scala 343:55]
  wire [31:0] _GEN_686 = _hit_T | writeBack ? _GEN_674 : _GEN_680; // @[dcache.scala 343:55]
  wire [127:0] _GEN_687 = _hit_T | writeBack ? _GEN_675 : _GEN_681; // @[dcache.scala 343:55]
  wire [2:0] _GEN_688 = _hit_T | writeBack ? _GEN_676 : _GEN_683; // @[dcache.scala 343:55]
  wire [3:0] _GEN_689 = _hit_T | writeBack ? _GEN_677 : _GEN_682; // @[dcache.scala 343:55]
  wire  _GEN_690 = _hit_T | writeBack ? 1'h0 : _T_43; // @[dcache.scala 157:25 343:55]
  wire [2:0] _GEN_691 = war_stall ? 3'h3 : _GEN_684; // @[dcache.scala 340:33 341:27]
  wire  _GEN_692 = war_stall ? 1'h0 : _GEN_685; // @[dcache.scala 161:25 340:33]
  wire [31:0] _GEN_693 = war_stall ? 32'h0 : _GEN_686; // @[dcache.scala 163:25 340:33]
  wire [127:0] _GEN_694 = war_stall ? 128'h0 : _GEN_687; // @[dcache.scala 165:25 340:33]
  wire [2:0] _GEN_695 = war_stall ? 3'h0 : _GEN_688; // @[dcache.scala 162:25 340:33]
  wire [3:0] _GEN_696 = war_stall ? 4'h0 : _GEN_689; // @[dcache.scala 164:25 340:33]
  wire  _GEN_697 = war_stall ? 1'h0 : _GEN_690; // @[dcache.scala 157:25 340:33]
  wire [2:0] _GEN_698 = wr_rdy ? _GEN_691 : 3'h3; // @[dcache.scala 334:23 339:31]
  wire  _GEN_699 = wr_rdy & _GEN_692; // @[dcache.scala 161:25 339:31]
  wire [31:0] _GEN_700 = wr_rdy ? _GEN_693 : 32'h0; // @[dcache.scala 163:25 339:31]
  wire [127:0] _GEN_701 = wr_rdy ? _GEN_694 : 128'h0; // @[dcache.scala 165:25 339:31]
  wire [2:0] _GEN_702 = wr_rdy ? _GEN_695 : 3'h0; // @[dcache.scala 162:25 339:31]
  wire [3:0] _GEN_703 = wr_rdy ? _GEN_696 : 4'h0; // @[dcache.scala 164:25 339:31]
  wire  _GEN_704 = wr_rdy & _GEN_697; // @[dcache.scala 157:25 339:31]
  wire [2:0] _GEN_705 = _T_6 & req_uncached ? 3'h4 : _GEN_698; // @[dcache.scala 336:42 337:25]
  wire  _GEN_706 = _T_6 & req_uncached ? 1'h0 : _GEN_699; // @[dcache.scala 161:25 336:42]
  wire [31:0] _GEN_707 = _T_6 & req_uncached ? 32'h0 : _GEN_700; // @[dcache.scala 163:25 336:42]
  wire [127:0] _GEN_708 = _T_6 & req_uncached ? 128'h0 : _GEN_701; // @[dcache.scala 165:25 336:42]
  wire [2:0] _GEN_709 = _T_6 & req_uncached ? 3'h0 : _GEN_702; // @[dcache.scala 162:25 336:42]
  wire [3:0] _GEN_710 = _T_6 & req_uncached ? 4'h0 : _GEN_703; // @[dcache.scala 164:25 336:42]
  wire  _GEN_711 = _T_6 & req_uncached ? 1'h0 : _GEN_704; // @[dcache.scala 157:25 336:42]
  wire  _rd_req_T_1 = _T_43 ? 1'h0 : 1'h1; // @[dcache.scala 368:39]
  wire [2:0] _rd_type_T_1 = req_uncached ? _wr_type_T : 3'h4; // @[dcache.scala 369:39]
  wire [31:0] _rd_addr_T_1 = {req_tag,req_set,4'h0}; // @[Cat.scala 33:92]
  wire [31:0] _rd_addr_T_2 = req_uncached ? _wr_addr_T_2 : _rd_addr_T_1; // @[dcache.scala 370:39]
  wire [2:0] _GEN_712 = rd_rdy ? 3'h5 : 3'h4; // @[dcache.scala 372:29 367:33 373:33]
  wire [2:0] _GEN_713 = _T_7 ? _GEN_712 : 3'h5; // @[dcache.scala 366:31 376:33]
  wire  _GEN_714 = _T_7 & _rd_req_T_1; // @[dcache.scala 158:25 366:31 368:33]
  wire [2:0] _GEN_715 = _T_7 ? _rd_type_T_1 : 3'h0; // @[dcache.scala 159:25 366:31 369:33]
  wire [31:0] _GEN_716 = _T_7 ? _rd_addr_T_2 : 32'h0; // @[dcache.scala 160:25 366:31 370:33]
  wire  _T_49 = _hit_T & _T_7; // @[dcache.scala 381:32]
  wire [1:0] _wr_cnt_T_1 = wr_cnt + 2'h1; // @[dcache.scala 385:71]
  wire  _GEN_12727 = 2'h0 == wr_cnt; // @[dcache.scala 149:33 386:{61,61}]
  wire [31:0] _GEN_717 = _GEN_11958 & 2'h0 == wr_cnt ? ret_data : 32'h0; // @[dcache.scala 149:33 386:{61,61}]
  wire  _GEN_12729 = 2'h1 == wr_cnt; // @[dcache.scala 149:33 386:{61,61}]
  wire [31:0] _GEN_718 = _GEN_11958 & 2'h1 == wr_cnt ? ret_data : 32'h0; // @[dcache.scala 149:33 386:{61,61}]
  wire  _GEN_12731 = 2'h2 == wr_cnt; // @[dcache.scala 149:33 386:{61,61}]
  wire [31:0] _GEN_719 = _GEN_11958 & 2'h2 == wr_cnt ? ret_data : 32'h0; // @[dcache.scala 149:33 386:{61,61}]
  wire  _GEN_12733 = 2'h3 == wr_cnt; // @[dcache.scala 149:33 386:{61,61}]
  wire [31:0] _GEN_720 = _GEN_11958 & 2'h3 == wr_cnt ? ret_data : 32'h0; // @[dcache.scala 149:33 386:{61,61}]
  wire [31:0] _GEN_721 = refillIDX_r & 2'h0 == wr_cnt ? ret_data : 32'h0; // @[dcache.scala 149:33 386:{61,61}]
  wire [31:0] _GEN_722 = refillIDX_r & 2'h1 == wr_cnt ? ret_data : 32'h0; // @[dcache.scala 149:33 386:{61,61}]
  wire [31:0] _GEN_723 = refillIDX_r & 2'h2 == wr_cnt ? ret_data : 32'h0; // @[dcache.scala 149:33 386:{61,61}]
  wire [31:0] _GEN_724 = refillIDX_r & 2'h3 == wr_cnt ? ret_data : 32'h0; // @[dcache.scala 149:33 386:{61,61}]
  wire [3:0] _GEN_725 = _GEN_11958 & _GEN_12727 ? 4'hf : 4'h0; // @[dcache.scala 150:33 387:{61,61}]
  wire [3:0] _GEN_726 = _GEN_11958 & _GEN_12729 ? 4'hf : 4'h0; // @[dcache.scala 150:33 387:{61,61}]
  wire [3:0] _GEN_727 = _GEN_11958 & _GEN_12731 ? 4'hf : 4'h0; // @[dcache.scala 150:33 387:{61,61}]
  wire [3:0] _GEN_728 = _GEN_11958 & _GEN_12733 ? 4'hf : 4'h0; // @[dcache.scala 150:33 387:{61,61}]
  wire [3:0] _GEN_729 = refillIDX_r & _GEN_12727 ? 4'hf : 4'h0; // @[dcache.scala 150:33 387:{61,61}]
  wire [3:0] _GEN_730 = refillIDX_r & _GEN_12729 ? 4'hf : 4'h0; // @[dcache.scala 150:33 387:{61,61}]
  wire [3:0] _GEN_731 = refillIDX_r & _GEN_12731 ? 4'hf : 4'h0; // @[dcache.scala 150:33 387:{61,61}]
  wire [3:0] _GEN_732 = refillIDX_r & _GEN_12733 ? 4'hf : 4'h0; // @[dcache.scala 150:33 387:{61,61}]
  wire  _GEN_733 = _GEN_11958 & _GEN_12468 ? 1'h0 : dirty_0_0; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_734 = _GEN_11958 & _GEN_11959 ? 1'h0 : dirty_0_1; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_735 = _GEN_11958 & _GEN_11961 ? 1'h0 : dirty_0_2; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_736 = _GEN_11958 & _GEN_11963 ? 1'h0 : dirty_0_3; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_737 = _GEN_11958 & _GEN_11965 ? 1'h0 : dirty_0_4; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_738 = _GEN_11958 & _GEN_11967 ? 1'h0 : dirty_0_5; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_739 = _GEN_11958 & _GEN_11969 ? 1'h0 : dirty_0_6; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_740 = _GEN_11958 & _GEN_11971 ? 1'h0 : dirty_0_7; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_741 = _GEN_11958 & _GEN_11973 ? 1'h0 : dirty_0_8; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_742 = _GEN_11958 & _GEN_11975 ? 1'h0 : dirty_0_9; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_743 = _GEN_11958 & _GEN_11977 ? 1'h0 : dirty_0_10; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_744 = _GEN_11958 & _GEN_11979 ? 1'h0 : dirty_0_11; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_745 = _GEN_11958 & _GEN_11981 ? 1'h0 : dirty_0_12; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_746 = _GEN_11958 & _GEN_11983 ? 1'h0 : dirty_0_13; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_747 = _GEN_11958 & _GEN_11985 ? 1'h0 : dirty_0_14; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_748 = _GEN_11958 & _GEN_11987 ? 1'h0 : dirty_0_15; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_749 = _GEN_11958 & _GEN_11989 ? 1'h0 : dirty_0_16; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_750 = _GEN_11958 & _GEN_11991 ? 1'h0 : dirty_0_17; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_751 = _GEN_11958 & _GEN_11993 ? 1'h0 : dirty_0_18; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_752 = _GEN_11958 & _GEN_11995 ? 1'h0 : dirty_0_19; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_753 = _GEN_11958 & _GEN_11997 ? 1'h0 : dirty_0_20; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_754 = _GEN_11958 & _GEN_11999 ? 1'h0 : dirty_0_21; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_755 = _GEN_11958 & _GEN_12001 ? 1'h0 : dirty_0_22; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_756 = _GEN_11958 & _GEN_12003 ? 1'h0 : dirty_0_23; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_757 = _GEN_11958 & _GEN_12005 ? 1'h0 : dirty_0_24; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_758 = _GEN_11958 & _GEN_12007 ? 1'h0 : dirty_0_25; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_759 = _GEN_11958 & _GEN_12009 ? 1'h0 : dirty_0_26; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_760 = _GEN_11958 & _GEN_12011 ? 1'h0 : dirty_0_27; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_761 = _GEN_11958 & _GEN_12013 ? 1'h0 : dirty_0_28; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_762 = _GEN_11958 & _GEN_12015 ? 1'h0 : dirty_0_29; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_763 = _GEN_11958 & _GEN_12017 ? 1'h0 : dirty_0_30; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_764 = _GEN_11958 & _GEN_12019 ? 1'h0 : dirty_0_31; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_765 = _GEN_11958 & _GEN_12021 ? 1'h0 : dirty_0_32; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_766 = _GEN_11958 & _GEN_12023 ? 1'h0 : dirty_0_33; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_767 = _GEN_11958 & _GEN_12025 ? 1'h0 : dirty_0_34; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_768 = _GEN_11958 & _GEN_12027 ? 1'h0 : dirty_0_35; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_769 = _GEN_11958 & _GEN_12029 ? 1'h0 : dirty_0_36; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_770 = _GEN_11958 & _GEN_12031 ? 1'h0 : dirty_0_37; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_771 = _GEN_11958 & _GEN_12033 ? 1'h0 : dirty_0_38; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_772 = _GEN_11958 & _GEN_12035 ? 1'h0 : dirty_0_39; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_773 = _GEN_11958 & _GEN_12037 ? 1'h0 : dirty_0_40; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_774 = _GEN_11958 & _GEN_12039 ? 1'h0 : dirty_0_41; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_775 = _GEN_11958 & _GEN_12041 ? 1'h0 : dirty_0_42; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_776 = _GEN_11958 & _GEN_12043 ? 1'h0 : dirty_0_43; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_777 = _GEN_11958 & _GEN_12045 ? 1'h0 : dirty_0_44; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_778 = _GEN_11958 & _GEN_12047 ? 1'h0 : dirty_0_45; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_779 = _GEN_11958 & _GEN_12049 ? 1'h0 : dirty_0_46; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_780 = _GEN_11958 & _GEN_12051 ? 1'h0 : dirty_0_47; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_781 = _GEN_11958 & _GEN_12053 ? 1'h0 : dirty_0_48; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_782 = _GEN_11958 & _GEN_12055 ? 1'h0 : dirty_0_49; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_783 = _GEN_11958 & _GEN_12057 ? 1'h0 : dirty_0_50; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_784 = _GEN_11958 & _GEN_12059 ? 1'h0 : dirty_0_51; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_785 = _GEN_11958 & _GEN_12061 ? 1'h0 : dirty_0_52; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_786 = _GEN_11958 & _GEN_12063 ? 1'h0 : dirty_0_53; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_787 = _GEN_11958 & _GEN_12065 ? 1'h0 : dirty_0_54; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_788 = _GEN_11958 & _GEN_12067 ? 1'h0 : dirty_0_55; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_789 = _GEN_11958 & _GEN_12069 ? 1'h0 : dirty_0_56; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_790 = _GEN_11958 & _GEN_12071 ? 1'h0 : dirty_0_57; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_791 = _GEN_11958 & _GEN_12073 ? 1'h0 : dirty_0_58; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_792 = _GEN_11958 & _GEN_12075 ? 1'h0 : dirty_0_59; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_793 = _GEN_11958 & _GEN_12077 ? 1'h0 : dirty_0_60; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_794 = _GEN_11958 & _GEN_12079 ? 1'h0 : dirty_0_61; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_795 = _GEN_11958 & _GEN_12081 ? 1'h0 : dirty_0_62; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_796 = _GEN_11958 & _GEN_12083 ? 1'h0 : dirty_0_63; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_797 = _GEN_11958 & _GEN_12085 ? 1'h0 : dirty_0_64; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_798 = _GEN_11958 & _GEN_12087 ? 1'h0 : dirty_0_65; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_799 = _GEN_11958 & _GEN_12089 ? 1'h0 : dirty_0_66; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_800 = _GEN_11958 & _GEN_12091 ? 1'h0 : dirty_0_67; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_801 = _GEN_11958 & _GEN_12093 ? 1'h0 : dirty_0_68; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_802 = _GEN_11958 & _GEN_12095 ? 1'h0 : dirty_0_69; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_803 = _GEN_11958 & _GEN_12097 ? 1'h0 : dirty_0_70; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_804 = _GEN_11958 & _GEN_12099 ? 1'h0 : dirty_0_71; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_805 = _GEN_11958 & _GEN_12101 ? 1'h0 : dirty_0_72; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_806 = _GEN_11958 & _GEN_12103 ? 1'h0 : dirty_0_73; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_807 = _GEN_11958 & _GEN_12105 ? 1'h0 : dirty_0_74; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_808 = _GEN_11958 & _GEN_12107 ? 1'h0 : dirty_0_75; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_809 = _GEN_11958 & _GEN_12109 ? 1'h0 : dirty_0_76; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_810 = _GEN_11958 & _GEN_12111 ? 1'h0 : dirty_0_77; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_811 = _GEN_11958 & _GEN_12113 ? 1'h0 : dirty_0_78; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_812 = _GEN_11958 & _GEN_12115 ? 1'h0 : dirty_0_79; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_813 = _GEN_11958 & _GEN_12117 ? 1'h0 : dirty_0_80; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_814 = _GEN_11958 & _GEN_12119 ? 1'h0 : dirty_0_81; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_815 = _GEN_11958 & _GEN_12121 ? 1'h0 : dirty_0_82; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_816 = _GEN_11958 & _GEN_12123 ? 1'h0 : dirty_0_83; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_817 = _GEN_11958 & _GEN_12125 ? 1'h0 : dirty_0_84; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_818 = _GEN_11958 & _GEN_12127 ? 1'h0 : dirty_0_85; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_819 = _GEN_11958 & _GEN_12129 ? 1'h0 : dirty_0_86; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_820 = _GEN_11958 & _GEN_12131 ? 1'h0 : dirty_0_87; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_821 = _GEN_11958 & _GEN_12133 ? 1'h0 : dirty_0_88; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_822 = _GEN_11958 & _GEN_12135 ? 1'h0 : dirty_0_89; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_823 = _GEN_11958 & _GEN_12137 ? 1'h0 : dirty_0_90; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_824 = _GEN_11958 & _GEN_12139 ? 1'h0 : dirty_0_91; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_825 = _GEN_11958 & _GEN_12141 ? 1'h0 : dirty_0_92; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_826 = _GEN_11958 & _GEN_12143 ? 1'h0 : dirty_0_93; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_827 = _GEN_11958 & _GEN_12145 ? 1'h0 : dirty_0_94; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_828 = _GEN_11958 & _GEN_12147 ? 1'h0 : dirty_0_95; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_829 = _GEN_11958 & _GEN_12149 ? 1'h0 : dirty_0_96; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_830 = _GEN_11958 & _GEN_12151 ? 1'h0 : dirty_0_97; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_831 = _GEN_11958 & _GEN_12153 ? 1'h0 : dirty_0_98; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_832 = _GEN_11958 & _GEN_12155 ? 1'h0 : dirty_0_99; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_833 = _GEN_11958 & _GEN_12157 ? 1'h0 : dirty_0_100; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_834 = _GEN_11958 & _GEN_12159 ? 1'h0 : dirty_0_101; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_835 = _GEN_11958 & _GEN_12161 ? 1'h0 : dirty_0_102; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_836 = _GEN_11958 & _GEN_12163 ? 1'h0 : dirty_0_103; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_837 = _GEN_11958 & _GEN_12165 ? 1'h0 : dirty_0_104; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_838 = _GEN_11958 & _GEN_12167 ? 1'h0 : dirty_0_105; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_839 = _GEN_11958 & _GEN_12169 ? 1'h0 : dirty_0_106; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_840 = _GEN_11958 & _GEN_12171 ? 1'h0 : dirty_0_107; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_841 = _GEN_11958 & _GEN_12173 ? 1'h0 : dirty_0_108; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_842 = _GEN_11958 & _GEN_12175 ? 1'h0 : dirty_0_109; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_843 = _GEN_11958 & _GEN_12177 ? 1'h0 : dirty_0_110; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_844 = _GEN_11958 & _GEN_12179 ? 1'h0 : dirty_0_111; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_845 = _GEN_11958 & _GEN_12181 ? 1'h0 : dirty_0_112; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_846 = _GEN_11958 & _GEN_12183 ? 1'h0 : dirty_0_113; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_847 = _GEN_11958 & _GEN_12185 ? 1'h0 : dirty_0_114; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_848 = _GEN_11958 & _GEN_12187 ? 1'h0 : dirty_0_115; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_849 = _GEN_11958 & _GEN_12189 ? 1'h0 : dirty_0_116; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_850 = _GEN_11958 & _GEN_12191 ? 1'h0 : dirty_0_117; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_851 = _GEN_11958 & _GEN_12193 ? 1'h0 : dirty_0_118; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_852 = _GEN_11958 & _GEN_12195 ? 1'h0 : dirty_0_119; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_853 = _GEN_11958 & _GEN_12197 ? 1'h0 : dirty_0_120; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_854 = _GEN_11958 & _GEN_12199 ? 1'h0 : dirty_0_121; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_855 = _GEN_11958 & _GEN_12201 ? 1'h0 : dirty_0_122; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_856 = _GEN_11958 & _GEN_12203 ? 1'h0 : dirty_0_123; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_857 = _GEN_11958 & _GEN_12205 ? 1'h0 : dirty_0_124; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_858 = _GEN_11958 & _GEN_12207 ? 1'h0 : dirty_0_125; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_859 = _GEN_11958 & _GEN_12209 ? 1'h0 : dirty_0_126; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_860 = _GEN_11958 & _GEN_12211 ? 1'h0 : dirty_0_127; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_861 = _GEN_11958 & _GEN_12213 ? 1'h0 : dirty_0_128; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_862 = _GEN_11958 & _GEN_12215 ? 1'h0 : dirty_0_129; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_863 = _GEN_11958 & _GEN_12217 ? 1'h0 : dirty_0_130; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_864 = _GEN_11958 & _GEN_12219 ? 1'h0 : dirty_0_131; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_865 = _GEN_11958 & _GEN_12221 ? 1'h0 : dirty_0_132; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_866 = _GEN_11958 & _GEN_12223 ? 1'h0 : dirty_0_133; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_867 = _GEN_11958 & _GEN_12225 ? 1'h0 : dirty_0_134; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_868 = _GEN_11958 & _GEN_12227 ? 1'h0 : dirty_0_135; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_869 = _GEN_11958 & _GEN_12229 ? 1'h0 : dirty_0_136; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_870 = _GEN_11958 & _GEN_12231 ? 1'h0 : dirty_0_137; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_871 = _GEN_11958 & _GEN_12233 ? 1'h0 : dirty_0_138; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_872 = _GEN_11958 & _GEN_12235 ? 1'h0 : dirty_0_139; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_873 = _GEN_11958 & _GEN_12237 ? 1'h0 : dirty_0_140; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_874 = _GEN_11958 & _GEN_12239 ? 1'h0 : dirty_0_141; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_875 = _GEN_11958 & _GEN_12241 ? 1'h0 : dirty_0_142; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_876 = _GEN_11958 & _GEN_12243 ? 1'h0 : dirty_0_143; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_877 = _GEN_11958 & _GEN_12245 ? 1'h0 : dirty_0_144; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_878 = _GEN_11958 & _GEN_12247 ? 1'h0 : dirty_0_145; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_879 = _GEN_11958 & _GEN_12249 ? 1'h0 : dirty_0_146; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_880 = _GEN_11958 & _GEN_12251 ? 1'h0 : dirty_0_147; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_881 = _GEN_11958 & _GEN_12253 ? 1'h0 : dirty_0_148; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_882 = _GEN_11958 & _GEN_12255 ? 1'h0 : dirty_0_149; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_883 = _GEN_11958 & _GEN_12257 ? 1'h0 : dirty_0_150; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_884 = _GEN_11958 & _GEN_12259 ? 1'h0 : dirty_0_151; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_885 = _GEN_11958 & _GEN_12261 ? 1'h0 : dirty_0_152; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_886 = _GEN_11958 & _GEN_12263 ? 1'h0 : dirty_0_153; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_887 = _GEN_11958 & _GEN_12265 ? 1'h0 : dirty_0_154; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_888 = _GEN_11958 & _GEN_12267 ? 1'h0 : dirty_0_155; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_889 = _GEN_11958 & _GEN_12269 ? 1'h0 : dirty_0_156; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_890 = _GEN_11958 & _GEN_12271 ? 1'h0 : dirty_0_157; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_891 = _GEN_11958 & _GEN_12273 ? 1'h0 : dirty_0_158; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_892 = _GEN_11958 & _GEN_12275 ? 1'h0 : dirty_0_159; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_893 = _GEN_11958 & _GEN_12277 ? 1'h0 : dirty_0_160; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_894 = _GEN_11958 & _GEN_12279 ? 1'h0 : dirty_0_161; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_895 = _GEN_11958 & _GEN_12281 ? 1'h0 : dirty_0_162; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_896 = _GEN_11958 & _GEN_12283 ? 1'h0 : dirty_0_163; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_897 = _GEN_11958 & _GEN_12285 ? 1'h0 : dirty_0_164; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_898 = _GEN_11958 & _GEN_12287 ? 1'h0 : dirty_0_165; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_899 = _GEN_11958 & _GEN_12289 ? 1'h0 : dirty_0_166; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_900 = _GEN_11958 & _GEN_12291 ? 1'h0 : dirty_0_167; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_901 = _GEN_11958 & _GEN_12293 ? 1'h0 : dirty_0_168; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_902 = _GEN_11958 & _GEN_12295 ? 1'h0 : dirty_0_169; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_903 = _GEN_11958 & _GEN_12297 ? 1'h0 : dirty_0_170; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_904 = _GEN_11958 & _GEN_12299 ? 1'h0 : dirty_0_171; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_905 = _GEN_11958 & _GEN_12301 ? 1'h0 : dirty_0_172; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_906 = _GEN_11958 & _GEN_12303 ? 1'h0 : dirty_0_173; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_907 = _GEN_11958 & _GEN_12305 ? 1'h0 : dirty_0_174; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_908 = _GEN_11958 & _GEN_12307 ? 1'h0 : dirty_0_175; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_909 = _GEN_11958 & _GEN_12309 ? 1'h0 : dirty_0_176; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_910 = _GEN_11958 & _GEN_12311 ? 1'h0 : dirty_0_177; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_911 = _GEN_11958 & _GEN_12313 ? 1'h0 : dirty_0_178; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_912 = _GEN_11958 & _GEN_12315 ? 1'h0 : dirty_0_179; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_913 = _GEN_11958 & _GEN_12317 ? 1'h0 : dirty_0_180; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_914 = _GEN_11958 & _GEN_12319 ? 1'h0 : dirty_0_181; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_915 = _GEN_11958 & _GEN_12321 ? 1'h0 : dirty_0_182; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_916 = _GEN_11958 & _GEN_12323 ? 1'h0 : dirty_0_183; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_917 = _GEN_11958 & _GEN_12325 ? 1'h0 : dirty_0_184; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_918 = _GEN_11958 & _GEN_12327 ? 1'h0 : dirty_0_185; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_919 = _GEN_11958 & _GEN_12329 ? 1'h0 : dirty_0_186; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_920 = _GEN_11958 & _GEN_12331 ? 1'h0 : dirty_0_187; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_921 = _GEN_11958 & _GEN_12333 ? 1'h0 : dirty_0_188; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_922 = _GEN_11958 & _GEN_12335 ? 1'h0 : dirty_0_189; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_923 = _GEN_11958 & _GEN_12337 ? 1'h0 : dirty_0_190; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_924 = _GEN_11958 & _GEN_12339 ? 1'h0 : dirty_0_191; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_925 = _GEN_11958 & _GEN_12341 ? 1'h0 : dirty_0_192; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_926 = _GEN_11958 & _GEN_12343 ? 1'h0 : dirty_0_193; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_927 = _GEN_11958 & _GEN_12345 ? 1'h0 : dirty_0_194; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_928 = _GEN_11958 & _GEN_12347 ? 1'h0 : dirty_0_195; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_929 = _GEN_11958 & _GEN_12349 ? 1'h0 : dirty_0_196; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_930 = _GEN_11958 & _GEN_12351 ? 1'h0 : dirty_0_197; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_931 = _GEN_11958 & _GEN_12353 ? 1'h0 : dirty_0_198; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_932 = _GEN_11958 & _GEN_12355 ? 1'h0 : dirty_0_199; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_933 = _GEN_11958 & _GEN_12357 ? 1'h0 : dirty_0_200; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_934 = _GEN_11958 & _GEN_12359 ? 1'h0 : dirty_0_201; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_935 = _GEN_11958 & _GEN_12361 ? 1'h0 : dirty_0_202; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_936 = _GEN_11958 & _GEN_12363 ? 1'h0 : dirty_0_203; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_937 = _GEN_11958 & _GEN_12365 ? 1'h0 : dirty_0_204; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_938 = _GEN_11958 & _GEN_12367 ? 1'h0 : dirty_0_205; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_939 = _GEN_11958 & _GEN_12369 ? 1'h0 : dirty_0_206; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_940 = _GEN_11958 & _GEN_12371 ? 1'h0 : dirty_0_207; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_941 = _GEN_11958 & _GEN_12373 ? 1'h0 : dirty_0_208; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_942 = _GEN_11958 & _GEN_12375 ? 1'h0 : dirty_0_209; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_943 = _GEN_11958 & _GEN_12377 ? 1'h0 : dirty_0_210; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_944 = _GEN_11958 & _GEN_12379 ? 1'h0 : dirty_0_211; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_945 = _GEN_11958 & _GEN_12381 ? 1'h0 : dirty_0_212; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_946 = _GEN_11958 & _GEN_12383 ? 1'h0 : dirty_0_213; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_947 = _GEN_11958 & _GEN_12385 ? 1'h0 : dirty_0_214; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_948 = _GEN_11958 & _GEN_12387 ? 1'h0 : dirty_0_215; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_949 = _GEN_11958 & _GEN_12389 ? 1'h0 : dirty_0_216; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_950 = _GEN_11958 & _GEN_12391 ? 1'h0 : dirty_0_217; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_951 = _GEN_11958 & _GEN_12393 ? 1'h0 : dirty_0_218; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_952 = _GEN_11958 & _GEN_12395 ? 1'h0 : dirty_0_219; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_953 = _GEN_11958 & _GEN_12397 ? 1'h0 : dirty_0_220; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_954 = _GEN_11958 & _GEN_12399 ? 1'h0 : dirty_0_221; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_955 = _GEN_11958 & _GEN_12401 ? 1'h0 : dirty_0_222; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_956 = _GEN_11958 & _GEN_12403 ? 1'h0 : dirty_0_223; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_957 = _GEN_11958 & _GEN_12405 ? 1'h0 : dirty_0_224; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_958 = _GEN_11958 & _GEN_12407 ? 1'h0 : dirty_0_225; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_959 = _GEN_11958 & _GEN_12409 ? 1'h0 : dirty_0_226; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_960 = _GEN_11958 & _GEN_12411 ? 1'h0 : dirty_0_227; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_961 = _GEN_11958 & _GEN_12413 ? 1'h0 : dirty_0_228; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_962 = _GEN_11958 & _GEN_12415 ? 1'h0 : dirty_0_229; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_963 = _GEN_11958 & _GEN_12417 ? 1'h0 : dirty_0_230; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_964 = _GEN_11958 & _GEN_12419 ? 1'h0 : dirty_0_231; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_965 = _GEN_11958 & _GEN_12421 ? 1'h0 : dirty_0_232; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_966 = _GEN_11958 & _GEN_12423 ? 1'h0 : dirty_0_233; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_967 = _GEN_11958 & _GEN_12425 ? 1'h0 : dirty_0_234; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_968 = _GEN_11958 & _GEN_12427 ? 1'h0 : dirty_0_235; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_969 = _GEN_11958 & _GEN_12429 ? 1'h0 : dirty_0_236; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_970 = _GEN_11958 & _GEN_12431 ? 1'h0 : dirty_0_237; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_971 = _GEN_11958 & _GEN_12433 ? 1'h0 : dirty_0_238; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_972 = _GEN_11958 & _GEN_12435 ? 1'h0 : dirty_0_239; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_973 = _GEN_11958 & _GEN_12437 ? 1'h0 : dirty_0_240; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_974 = _GEN_11958 & _GEN_12439 ? 1'h0 : dirty_0_241; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_975 = _GEN_11958 & _GEN_12441 ? 1'h0 : dirty_0_242; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_976 = _GEN_11958 & _GEN_12443 ? 1'h0 : dirty_0_243; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_977 = _GEN_11958 & _GEN_12445 ? 1'h0 : dirty_0_244; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_978 = _GEN_11958 & _GEN_12447 ? 1'h0 : dirty_0_245; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_979 = _GEN_11958 & _GEN_12449 ? 1'h0 : dirty_0_246; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_980 = _GEN_11958 & _GEN_12451 ? 1'h0 : dirty_0_247; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_981 = _GEN_11958 & _GEN_12453 ? 1'h0 : dirty_0_248; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_982 = _GEN_11958 & _GEN_12455 ? 1'h0 : dirty_0_249; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_983 = _GEN_11958 & _GEN_12457 ? 1'h0 : dirty_0_250; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_984 = _GEN_11958 & _GEN_12459 ? 1'h0 : dirty_0_251; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_985 = _GEN_11958 & _GEN_12461 ? 1'h0 : dirty_0_252; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_986 = _GEN_11958 & _GEN_12463 ? 1'h0 : dirty_0_253; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_987 = _GEN_11958 & _GEN_12465 ? 1'h0 : dirty_0_254; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_988 = _GEN_11958 & _GEN_12467 ? 1'h0 : dirty_0_255; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_989 = refillIDX_r & _GEN_12468 ? 1'h0 : dirty_1_0; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_990 = refillIDX_r & _GEN_11959 ? 1'h0 : dirty_1_1; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_991 = refillIDX_r & _GEN_11961 ? 1'h0 : dirty_1_2; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_992 = refillIDX_r & _GEN_11963 ? 1'h0 : dirty_1_3; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_993 = refillIDX_r & _GEN_11965 ? 1'h0 : dirty_1_4; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_994 = refillIDX_r & _GEN_11967 ? 1'h0 : dirty_1_5; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_995 = refillIDX_r & _GEN_11969 ? 1'h0 : dirty_1_6; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_996 = refillIDX_r & _GEN_11971 ? 1'h0 : dirty_1_7; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_997 = refillIDX_r & _GEN_11973 ? 1'h0 : dirty_1_8; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_998 = refillIDX_r & _GEN_11975 ? 1'h0 : dirty_1_9; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_999 = refillIDX_r & _GEN_11977 ? 1'h0 : dirty_1_10; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1000 = refillIDX_r & _GEN_11979 ? 1'h0 : dirty_1_11; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1001 = refillIDX_r & _GEN_11981 ? 1'h0 : dirty_1_12; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1002 = refillIDX_r & _GEN_11983 ? 1'h0 : dirty_1_13; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1003 = refillIDX_r & _GEN_11985 ? 1'h0 : dirty_1_14; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1004 = refillIDX_r & _GEN_11987 ? 1'h0 : dirty_1_15; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1005 = refillIDX_r & _GEN_11989 ? 1'h0 : dirty_1_16; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1006 = refillIDX_r & _GEN_11991 ? 1'h0 : dirty_1_17; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1007 = refillIDX_r & _GEN_11993 ? 1'h0 : dirty_1_18; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1008 = refillIDX_r & _GEN_11995 ? 1'h0 : dirty_1_19; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1009 = refillIDX_r & _GEN_11997 ? 1'h0 : dirty_1_20; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1010 = refillIDX_r & _GEN_11999 ? 1'h0 : dirty_1_21; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1011 = refillIDX_r & _GEN_12001 ? 1'h0 : dirty_1_22; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1012 = refillIDX_r & _GEN_12003 ? 1'h0 : dirty_1_23; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1013 = refillIDX_r & _GEN_12005 ? 1'h0 : dirty_1_24; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1014 = refillIDX_r & _GEN_12007 ? 1'h0 : dirty_1_25; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1015 = refillIDX_r & _GEN_12009 ? 1'h0 : dirty_1_26; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1016 = refillIDX_r & _GEN_12011 ? 1'h0 : dirty_1_27; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1017 = refillIDX_r & _GEN_12013 ? 1'h0 : dirty_1_28; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1018 = refillIDX_r & _GEN_12015 ? 1'h0 : dirty_1_29; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1019 = refillIDX_r & _GEN_12017 ? 1'h0 : dirty_1_30; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1020 = refillIDX_r & _GEN_12019 ? 1'h0 : dirty_1_31; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1021 = refillIDX_r & _GEN_12021 ? 1'h0 : dirty_1_32; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1022 = refillIDX_r & _GEN_12023 ? 1'h0 : dirty_1_33; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1023 = refillIDX_r & _GEN_12025 ? 1'h0 : dirty_1_34; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1024 = refillIDX_r & _GEN_12027 ? 1'h0 : dirty_1_35; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1025 = refillIDX_r & _GEN_12029 ? 1'h0 : dirty_1_36; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1026 = refillIDX_r & _GEN_12031 ? 1'h0 : dirty_1_37; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1027 = refillIDX_r & _GEN_12033 ? 1'h0 : dirty_1_38; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1028 = refillIDX_r & _GEN_12035 ? 1'h0 : dirty_1_39; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1029 = refillIDX_r & _GEN_12037 ? 1'h0 : dirty_1_40; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1030 = refillIDX_r & _GEN_12039 ? 1'h0 : dirty_1_41; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1031 = refillIDX_r & _GEN_12041 ? 1'h0 : dirty_1_42; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1032 = refillIDX_r & _GEN_12043 ? 1'h0 : dirty_1_43; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1033 = refillIDX_r & _GEN_12045 ? 1'h0 : dirty_1_44; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1034 = refillIDX_r & _GEN_12047 ? 1'h0 : dirty_1_45; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1035 = refillIDX_r & _GEN_12049 ? 1'h0 : dirty_1_46; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1036 = refillIDX_r & _GEN_12051 ? 1'h0 : dirty_1_47; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1037 = refillIDX_r & _GEN_12053 ? 1'h0 : dirty_1_48; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1038 = refillIDX_r & _GEN_12055 ? 1'h0 : dirty_1_49; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1039 = refillIDX_r & _GEN_12057 ? 1'h0 : dirty_1_50; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1040 = refillIDX_r & _GEN_12059 ? 1'h0 : dirty_1_51; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1041 = refillIDX_r & _GEN_12061 ? 1'h0 : dirty_1_52; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1042 = refillIDX_r & _GEN_12063 ? 1'h0 : dirty_1_53; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1043 = refillIDX_r & _GEN_12065 ? 1'h0 : dirty_1_54; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1044 = refillIDX_r & _GEN_12067 ? 1'h0 : dirty_1_55; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1045 = refillIDX_r & _GEN_12069 ? 1'h0 : dirty_1_56; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1046 = refillIDX_r & _GEN_12071 ? 1'h0 : dirty_1_57; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1047 = refillIDX_r & _GEN_12073 ? 1'h0 : dirty_1_58; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1048 = refillIDX_r & _GEN_12075 ? 1'h0 : dirty_1_59; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1049 = refillIDX_r & _GEN_12077 ? 1'h0 : dirty_1_60; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1050 = refillIDX_r & _GEN_12079 ? 1'h0 : dirty_1_61; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1051 = refillIDX_r & _GEN_12081 ? 1'h0 : dirty_1_62; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1052 = refillIDX_r & _GEN_12083 ? 1'h0 : dirty_1_63; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1053 = refillIDX_r & _GEN_12085 ? 1'h0 : dirty_1_64; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1054 = refillIDX_r & _GEN_12087 ? 1'h0 : dirty_1_65; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1055 = refillIDX_r & _GEN_12089 ? 1'h0 : dirty_1_66; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1056 = refillIDX_r & _GEN_12091 ? 1'h0 : dirty_1_67; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1057 = refillIDX_r & _GEN_12093 ? 1'h0 : dirty_1_68; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1058 = refillIDX_r & _GEN_12095 ? 1'h0 : dirty_1_69; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1059 = refillIDX_r & _GEN_12097 ? 1'h0 : dirty_1_70; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1060 = refillIDX_r & _GEN_12099 ? 1'h0 : dirty_1_71; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1061 = refillIDX_r & _GEN_12101 ? 1'h0 : dirty_1_72; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1062 = refillIDX_r & _GEN_12103 ? 1'h0 : dirty_1_73; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1063 = refillIDX_r & _GEN_12105 ? 1'h0 : dirty_1_74; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1064 = refillIDX_r & _GEN_12107 ? 1'h0 : dirty_1_75; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1065 = refillIDX_r & _GEN_12109 ? 1'h0 : dirty_1_76; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1066 = refillIDX_r & _GEN_12111 ? 1'h0 : dirty_1_77; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1067 = refillIDX_r & _GEN_12113 ? 1'h0 : dirty_1_78; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1068 = refillIDX_r & _GEN_12115 ? 1'h0 : dirty_1_79; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1069 = refillIDX_r & _GEN_12117 ? 1'h0 : dirty_1_80; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1070 = refillIDX_r & _GEN_12119 ? 1'h0 : dirty_1_81; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1071 = refillIDX_r & _GEN_12121 ? 1'h0 : dirty_1_82; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1072 = refillIDX_r & _GEN_12123 ? 1'h0 : dirty_1_83; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1073 = refillIDX_r & _GEN_12125 ? 1'h0 : dirty_1_84; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1074 = refillIDX_r & _GEN_12127 ? 1'h0 : dirty_1_85; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1075 = refillIDX_r & _GEN_12129 ? 1'h0 : dirty_1_86; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1076 = refillIDX_r & _GEN_12131 ? 1'h0 : dirty_1_87; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1077 = refillIDX_r & _GEN_12133 ? 1'h0 : dirty_1_88; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1078 = refillIDX_r & _GEN_12135 ? 1'h0 : dirty_1_89; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1079 = refillIDX_r & _GEN_12137 ? 1'h0 : dirty_1_90; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1080 = refillIDX_r & _GEN_12139 ? 1'h0 : dirty_1_91; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1081 = refillIDX_r & _GEN_12141 ? 1'h0 : dirty_1_92; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1082 = refillIDX_r & _GEN_12143 ? 1'h0 : dirty_1_93; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1083 = refillIDX_r & _GEN_12145 ? 1'h0 : dirty_1_94; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1084 = refillIDX_r & _GEN_12147 ? 1'h0 : dirty_1_95; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1085 = refillIDX_r & _GEN_12149 ? 1'h0 : dirty_1_96; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1086 = refillIDX_r & _GEN_12151 ? 1'h0 : dirty_1_97; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1087 = refillIDX_r & _GEN_12153 ? 1'h0 : dirty_1_98; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1088 = refillIDX_r & _GEN_12155 ? 1'h0 : dirty_1_99; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1089 = refillIDX_r & _GEN_12157 ? 1'h0 : dirty_1_100; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1090 = refillIDX_r & _GEN_12159 ? 1'h0 : dirty_1_101; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1091 = refillIDX_r & _GEN_12161 ? 1'h0 : dirty_1_102; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1092 = refillIDX_r & _GEN_12163 ? 1'h0 : dirty_1_103; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1093 = refillIDX_r & _GEN_12165 ? 1'h0 : dirty_1_104; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1094 = refillIDX_r & _GEN_12167 ? 1'h0 : dirty_1_105; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1095 = refillIDX_r & _GEN_12169 ? 1'h0 : dirty_1_106; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1096 = refillIDX_r & _GEN_12171 ? 1'h0 : dirty_1_107; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1097 = refillIDX_r & _GEN_12173 ? 1'h0 : dirty_1_108; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1098 = refillIDX_r & _GEN_12175 ? 1'h0 : dirty_1_109; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1099 = refillIDX_r & _GEN_12177 ? 1'h0 : dirty_1_110; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1100 = refillIDX_r & _GEN_12179 ? 1'h0 : dirty_1_111; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1101 = refillIDX_r & _GEN_12181 ? 1'h0 : dirty_1_112; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1102 = refillIDX_r & _GEN_12183 ? 1'h0 : dirty_1_113; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1103 = refillIDX_r & _GEN_12185 ? 1'h0 : dirty_1_114; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1104 = refillIDX_r & _GEN_12187 ? 1'h0 : dirty_1_115; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1105 = refillIDX_r & _GEN_12189 ? 1'h0 : dirty_1_116; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1106 = refillIDX_r & _GEN_12191 ? 1'h0 : dirty_1_117; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1107 = refillIDX_r & _GEN_12193 ? 1'h0 : dirty_1_118; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1108 = refillIDX_r & _GEN_12195 ? 1'h0 : dirty_1_119; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1109 = refillIDX_r & _GEN_12197 ? 1'h0 : dirty_1_120; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1110 = refillIDX_r & _GEN_12199 ? 1'h0 : dirty_1_121; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1111 = refillIDX_r & _GEN_12201 ? 1'h0 : dirty_1_122; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1112 = refillIDX_r & _GEN_12203 ? 1'h0 : dirty_1_123; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1113 = refillIDX_r & _GEN_12205 ? 1'h0 : dirty_1_124; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1114 = refillIDX_r & _GEN_12207 ? 1'h0 : dirty_1_125; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1115 = refillIDX_r & _GEN_12209 ? 1'h0 : dirty_1_126; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1116 = refillIDX_r & _GEN_12211 ? 1'h0 : dirty_1_127; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1117 = refillIDX_r & _GEN_12213 ? 1'h0 : dirty_1_128; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1118 = refillIDX_r & _GEN_12215 ? 1'h0 : dirty_1_129; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1119 = refillIDX_r & _GEN_12217 ? 1'h0 : dirty_1_130; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1120 = refillIDX_r & _GEN_12219 ? 1'h0 : dirty_1_131; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1121 = refillIDX_r & _GEN_12221 ? 1'h0 : dirty_1_132; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1122 = refillIDX_r & _GEN_12223 ? 1'h0 : dirty_1_133; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1123 = refillIDX_r & _GEN_12225 ? 1'h0 : dirty_1_134; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1124 = refillIDX_r & _GEN_12227 ? 1'h0 : dirty_1_135; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1125 = refillIDX_r & _GEN_12229 ? 1'h0 : dirty_1_136; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1126 = refillIDX_r & _GEN_12231 ? 1'h0 : dirty_1_137; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1127 = refillIDX_r & _GEN_12233 ? 1'h0 : dirty_1_138; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1128 = refillIDX_r & _GEN_12235 ? 1'h0 : dirty_1_139; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1129 = refillIDX_r & _GEN_12237 ? 1'h0 : dirty_1_140; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1130 = refillIDX_r & _GEN_12239 ? 1'h0 : dirty_1_141; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1131 = refillIDX_r & _GEN_12241 ? 1'h0 : dirty_1_142; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1132 = refillIDX_r & _GEN_12243 ? 1'h0 : dirty_1_143; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1133 = refillIDX_r & _GEN_12245 ? 1'h0 : dirty_1_144; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1134 = refillIDX_r & _GEN_12247 ? 1'h0 : dirty_1_145; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1135 = refillIDX_r & _GEN_12249 ? 1'h0 : dirty_1_146; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1136 = refillIDX_r & _GEN_12251 ? 1'h0 : dirty_1_147; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1137 = refillIDX_r & _GEN_12253 ? 1'h0 : dirty_1_148; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1138 = refillIDX_r & _GEN_12255 ? 1'h0 : dirty_1_149; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1139 = refillIDX_r & _GEN_12257 ? 1'h0 : dirty_1_150; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1140 = refillIDX_r & _GEN_12259 ? 1'h0 : dirty_1_151; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1141 = refillIDX_r & _GEN_12261 ? 1'h0 : dirty_1_152; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1142 = refillIDX_r & _GEN_12263 ? 1'h0 : dirty_1_153; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1143 = refillIDX_r & _GEN_12265 ? 1'h0 : dirty_1_154; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1144 = refillIDX_r & _GEN_12267 ? 1'h0 : dirty_1_155; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1145 = refillIDX_r & _GEN_12269 ? 1'h0 : dirty_1_156; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1146 = refillIDX_r & _GEN_12271 ? 1'h0 : dirty_1_157; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1147 = refillIDX_r & _GEN_12273 ? 1'h0 : dirty_1_158; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1148 = refillIDX_r & _GEN_12275 ? 1'h0 : dirty_1_159; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1149 = refillIDX_r & _GEN_12277 ? 1'h0 : dirty_1_160; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1150 = refillIDX_r & _GEN_12279 ? 1'h0 : dirty_1_161; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1151 = refillIDX_r & _GEN_12281 ? 1'h0 : dirty_1_162; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1152 = refillIDX_r & _GEN_12283 ? 1'h0 : dirty_1_163; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1153 = refillIDX_r & _GEN_12285 ? 1'h0 : dirty_1_164; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1154 = refillIDX_r & _GEN_12287 ? 1'h0 : dirty_1_165; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1155 = refillIDX_r & _GEN_12289 ? 1'h0 : dirty_1_166; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1156 = refillIDX_r & _GEN_12291 ? 1'h0 : dirty_1_167; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1157 = refillIDX_r & _GEN_12293 ? 1'h0 : dirty_1_168; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1158 = refillIDX_r & _GEN_12295 ? 1'h0 : dirty_1_169; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1159 = refillIDX_r & _GEN_12297 ? 1'h0 : dirty_1_170; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1160 = refillIDX_r & _GEN_12299 ? 1'h0 : dirty_1_171; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1161 = refillIDX_r & _GEN_12301 ? 1'h0 : dirty_1_172; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1162 = refillIDX_r & _GEN_12303 ? 1'h0 : dirty_1_173; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1163 = refillIDX_r & _GEN_12305 ? 1'h0 : dirty_1_174; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1164 = refillIDX_r & _GEN_12307 ? 1'h0 : dirty_1_175; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1165 = refillIDX_r & _GEN_12309 ? 1'h0 : dirty_1_176; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1166 = refillIDX_r & _GEN_12311 ? 1'h0 : dirty_1_177; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1167 = refillIDX_r & _GEN_12313 ? 1'h0 : dirty_1_178; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1168 = refillIDX_r & _GEN_12315 ? 1'h0 : dirty_1_179; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1169 = refillIDX_r & _GEN_12317 ? 1'h0 : dirty_1_180; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1170 = refillIDX_r & _GEN_12319 ? 1'h0 : dirty_1_181; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1171 = refillIDX_r & _GEN_12321 ? 1'h0 : dirty_1_182; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1172 = refillIDX_r & _GEN_12323 ? 1'h0 : dirty_1_183; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1173 = refillIDX_r & _GEN_12325 ? 1'h0 : dirty_1_184; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1174 = refillIDX_r & _GEN_12327 ? 1'h0 : dirty_1_185; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1175 = refillIDX_r & _GEN_12329 ? 1'h0 : dirty_1_186; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1176 = refillIDX_r & _GEN_12331 ? 1'h0 : dirty_1_187; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1177 = refillIDX_r & _GEN_12333 ? 1'h0 : dirty_1_188; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1178 = refillIDX_r & _GEN_12335 ? 1'h0 : dirty_1_189; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1179 = refillIDX_r & _GEN_12337 ? 1'h0 : dirty_1_190; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1180 = refillIDX_r & _GEN_12339 ? 1'h0 : dirty_1_191; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1181 = refillIDX_r & _GEN_12341 ? 1'h0 : dirty_1_192; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1182 = refillIDX_r & _GEN_12343 ? 1'h0 : dirty_1_193; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1183 = refillIDX_r & _GEN_12345 ? 1'h0 : dirty_1_194; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1184 = refillIDX_r & _GEN_12347 ? 1'h0 : dirty_1_195; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1185 = refillIDX_r & _GEN_12349 ? 1'h0 : dirty_1_196; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1186 = refillIDX_r & _GEN_12351 ? 1'h0 : dirty_1_197; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1187 = refillIDX_r & _GEN_12353 ? 1'h0 : dirty_1_198; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1188 = refillIDX_r & _GEN_12355 ? 1'h0 : dirty_1_199; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1189 = refillIDX_r & _GEN_12357 ? 1'h0 : dirty_1_200; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1190 = refillIDX_r & _GEN_12359 ? 1'h0 : dirty_1_201; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1191 = refillIDX_r & _GEN_12361 ? 1'h0 : dirty_1_202; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1192 = refillIDX_r & _GEN_12363 ? 1'h0 : dirty_1_203; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1193 = refillIDX_r & _GEN_12365 ? 1'h0 : dirty_1_204; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1194 = refillIDX_r & _GEN_12367 ? 1'h0 : dirty_1_205; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1195 = refillIDX_r & _GEN_12369 ? 1'h0 : dirty_1_206; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1196 = refillIDX_r & _GEN_12371 ? 1'h0 : dirty_1_207; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1197 = refillIDX_r & _GEN_12373 ? 1'h0 : dirty_1_208; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1198 = refillIDX_r & _GEN_12375 ? 1'h0 : dirty_1_209; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1199 = refillIDX_r & _GEN_12377 ? 1'h0 : dirty_1_210; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1200 = refillIDX_r & _GEN_12379 ? 1'h0 : dirty_1_211; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1201 = refillIDX_r & _GEN_12381 ? 1'h0 : dirty_1_212; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1202 = refillIDX_r & _GEN_12383 ? 1'h0 : dirty_1_213; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1203 = refillIDX_r & _GEN_12385 ? 1'h0 : dirty_1_214; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1204 = refillIDX_r & _GEN_12387 ? 1'h0 : dirty_1_215; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1205 = refillIDX_r & _GEN_12389 ? 1'h0 : dirty_1_216; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1206 = refillIDX_r & _GEN_12391 ? 1'h0 : dirty_1_217; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1207 = refillIDX_r & _GEN_12393 ? 1'h0 : dirty_1_218; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1208 = refillIDX_r & _GEN_12395 ? 1'h0 : dirty_1_219; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1209 = refillIDX_r & _GEN_12397 ? 1'h0 : dirty_1_220; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1210 = refillIDX_r & _GEN_12399 ? 1'h0 : dirty_1_221; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1211 = refillIDX_r & _GEN_12401 ? 1'h0 : dirty_1_222; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1212 = refillIDX_r & _GEN_12403 ? 1'h0 : dirty_1_223; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1213 = refillIDX_r & _GEN_12405 ? 1'h0 : dirty_1_224; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1214 = refillIDX_r & _GEN_12407 ? 1'h0 : dirty_1_225; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1215 = refillIDX_r & _GEN_12409 ? 1'h0 : dirty_1_226; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1216 = refillIDX_r & _GEN_12411 ? 1'h0 : dirty_1_227; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1217 = refillIDX_r & _GEN_12413 ? 1'h0 : dirty_1_228; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1218 = refillIDX_r & _GEN_12415 ? 1'h0 : dirty_1_229; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1219 = refillIDX_r & _GEN_12417 ? 1'h0 : dirty_1_230; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1220 = refillIDX_r & _GEN_12419 ? 1'h0 : dirty_1_231; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1221 = refillIDX_r & _GEN_12421 ? 1'h0 : dirty_1_232; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1222 = refillIDX_r & _GEN_12423 ? 1'h0 : dirty_1_233; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1223 = refillIDX_r & _GEN_12425 ? 1'h0 : dirty_1_234; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1224 = refillIDX_r & _GEN_12427 ? 1'h0 : dirty_1_235; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1225 = refillIDX_r & _GEN_12429 ? 1'h0 : dirty_1_236; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1226 = refillIDX_r & _GEN_12431 ? 1'h0 : dirty_1_237; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1227 = refillIDX_r & _GEN_12433 ? 1'h0 : dirty_1_238; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1228 = refillIDX_r & _GEN_12435 ? 1'h0 : dirty_1_239; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1229 = refillIDX_r & _GEN_12437 ? 1'h0 : dirty_1_240; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1230 = refillIDX_r & _GEN_12439 ? 1'h0 : dirty_1_241; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1231 = refillIDX_r & _GEN_12441 ? 1'h0 : dirty_1_242; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1232 = refillIDX_r & _GEN_12443 ? 1'h0 : dirty_1_243; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1233 = refillIDX_r & _GEN_12445 ? 1'h0 : dirty_1_244; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1234 = refillIDX_r & _GEN_12447 ? 1'h0 : dirty_1_245; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1235 = refillIDX_r & _GEN_12449 ? 1'h0 : dirty_1_246; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1236 = refillIDX_r & _GEN_12451 ? 1'h0 : dirty_1_247; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1237 = refillIDX_r & _GEN_12453 ? 1'h0 : dirty_1_248; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1238 = refillIDX_r & _GEN_12455 ? 1'h0 : dirty_1_249; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1239 = refillIDX_r & _GEN_12457 ? 1'h0 : dirty_1_250; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1240 = refillIDX_r & _GEN_12459 ? 1'h0 : dirty_1_251; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1241 = refillIDX_r & _GEN_12461 ? 1'h0 : dirty_1_252; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1242 = refillIDX_r & _GEN_12463 ? 1'h0 : dirty_1_253; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1243 = refillIDX_r & _GEN_12465 ? 1'h0 : dirty_1_254; // @[dcache.scala 113:28 391:{61,61}]
  wire  _GEN_1244 = refillIDX_r & _GEN_12467 ? 1'h0 : dirty_1_255; // @[dcache.scala 113:28 391:{61,61}]
  wire [20:0] _tagv_dina_T = {1'h1,req_tag}; // @[Cat.scala 33:92]
  wire [20:0] _GEN_1247 = ~refillIDX_r ? _tagv_dina_T : 21'h0; // @[dcache.scala 143:25 393:{61,61}]
  wire [20:0] _GEN_1248 = refillIDX_r ? _tagv_dina_T : 21'h0; // @[dcache.scala 143:25 393:{61,61}]
  wire [2:0] _GEN_1249 = ret_last ? 3'h1 : 3'h5; // @[dcache.scala 389:21 380:41 390:61]
  wire  _GEN_1250 = ret_last ? _GEN_733 : dirty_0_0; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1251 = ret_last ? _GEN_734 : dirty_0_1; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1252 = ret_last ? _GEN_735 : dirty_0_2; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1253 = ret_last ? _GEN_736 : dirty_0_3; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1254 = ret_last ? _GEN_737 : dirty_0_4; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1255 = ret_last ? _GEN_738 : dirty_0_5; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1256 = ret_last ? _GEN_739 : dirty_0_6; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1257 = ret_last ? _GEN_740 : dirty_0_7; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1258 = ret_last ? _GEN_741 : dirty_0_8; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1259 = ret_last ? _GEN_742 : dirty_0_9; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1260 = ret_last ? _GEN_743 : dirty_0_10; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1261 = ret_last ? _GEN_744 : dirty_0_11; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1262 = ret_last ? _GEN_745 : dirty_0_12; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1263 = ret_last ? _GEN_746 : dirty_0_13; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1264 = ret_last ? _GEN_747 : dirty_0_14; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1265 = ret_last ? _GEN_748 : dirty_0_15; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1266 = ret_last ? _GEN_749 : dirty_0_16; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1267 = ret_last ? _GEN_750 : dirty_0_17; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1268 = ret_last ? _GEN_751 : dirty_0_18; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1269 = ret_last ? _GEN_752 : dirty_0_19; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1270 = ret_last ? _GEN_753 : dirty_0_20; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1271 = ret_last ? _GEN_754 : dirty_0_21; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1272 = ret_last ? _GEN_755 : dirty_0_22; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1273 = ret_last ? _GEN_756 : dirty_0_23; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1274 = ret_last ? _GEN_757 : dirty_0_24; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1275 = ret_last ? _GEN_758 : dirty_0_25; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1276 = ret_last ? _GEN_759 : dirty_0_26; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1277 = ret_last ? _GEN_760 : dirty_0_27; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1278 = ret_last ? _GEN_761 : dirty_0_28; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1279 = ret_last ? _GEN_762 : dirty_0_29; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1280 = ret_last ? _GEN_763 : dirty_0_30; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1281 = ret_last ? _GEN_764 : dirty_0_31; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1282 = ret_last ? _GEN_765 : dirty_0_32; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1283 = ret_last ? _GEN_766 : dirty_0_33; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1284 = ret_last ? _GEN_767 : dirty_0_34; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1285 = ret_last ? _GEN_768 : dirty_0_35; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1286 = ret_last ? _GEN_769 : dirty_0_36; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1287 = ret_last ? _GEN_770 : dirty_0_37; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1288 = ret_last ? _GEN_771 : dirty_0_38; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1289 = ret_last ? _GEN_772 : dirty_0_39; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1290 = ret_last ? _GEN_773 : dirty_0_40; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1291 = ret_last ? _GEN_774 : dirty_0_41; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1292 = ret_last ? _GEN_775 : dirty_0_42; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1293 = ret_last ? _GEN_776 : dirty_0_43; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1294 = ret_last ? _GEN_777 : dirty_0_44; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1295 = ret_last ? _GEN_778 : dirty_0_45; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1296 = ret_last ? _GEN_779 : dirty_0_46; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1297 = ret_last ? _GEN_780 : dirty_0_47; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1298 = ret_last ? _GEN_781 : dirty_0_48; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1299 = ret_last ? _GEN_782 : dirty_0_49; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1300 = ret_last ? _GEN_783 : dirty_0_50; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1301 = ret_last ? _GEN_784 : dirty_0_51; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1302 = ret_last ? _GEN_785 : dirty_0_52; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1303 = ret_last ? _GEN_786 : dirty_0_53; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1304 = ret_last ? _GEN_787 : dirty_0_54; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1305 = ret_last ? _GEN_788 : dirty_0_55; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1306 = ret_last ? _GEN_789 : dirty_0_56; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1307 = ret_last ? _GEN_790 : dirty_0_57; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1308 = ret_last ? _GEN_791 : dirty_0_58; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1309 = ret_last ? _GEN_792 : dirty_0_59; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1310 = ret_last ? _GEN_793 : dirty_0_60; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1311 = ret_last ? _GEN_794 : dirty_0_61; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1312 = ret_last ? _GEN_795 : dirty_0_62; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1313 = ret_last ? _GEN_796 : dirty_0_63; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1314 = ret_last ? _GEN_797 : dirty_0_64; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1315 = ret_last ? _GEN_798 : dirty_0_65; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1316 = ret_last ? _GEN_799 : dirty_0_66; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1317 = ret_last ? _GEN_800 : dirty_0_67; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1318 = ret_last ? _GEN_801 : dirty_0_68; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1319 = ret_last ? _GEN_802 : dirty_0_69; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1320 = ret_last ? _GEN_803 : dirty_0_70; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1321 = ret_last ? _GEN_804 : dirty_0_71; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1322 = ret_last ? _GEN_805 : dirty_0_72; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1323 = ret_last ? _GEN_806 : dirty_0_73; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1324 = ret_last ? _GEN_807 : dirty_0_74; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1325 = ret_last ? _GEN_808 : dirty_0_75; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1326 = ret_last ? _GEN_809 : dirty_0_76; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1327 = ret_last ? _GEN_810 : dirty_0_77; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1328 = ret_last ? _GEN_811 : dirty_0_78; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1329 = ret_last ? _GEN_812 : dirty_0_79; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1330 = ret_last ? _GEN_813 : dirty_0_80; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1331 = ret_last ? _GEN_814 : dirty_0_81; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1332 = ret_last ? _GEN_815 : dirty_0_82; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1333 = ret_last ? _GEN_816 : dirty_0_83; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1334 = ret_last ? _GEN_817 : dirty_0_84; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1335 = ret_last ? _GEN_818 : dirty_0_85; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1336 = ret_last ? _GEN_819 : dirty_0_86; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1337 = ret_last ? _GEN_820 : dirty_0_87; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1338 = ret_last ? _GEN_821 : dirty_0_88; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1339 = ret_last ? _GEN_822 : dirty_0_89; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1340 = ret_last ? _GEN_823 : dirty_0_90; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1341 = ret_last ? _GEN_824 : dirty_0_91; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1342 = ret_last ? _GEN_825 : dirty_0_92; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1343 = ret_last ? _GEN_826 : dirty_0_93; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1344 = ret_last ? _GEN_827 : dirty_0_94; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1345 = ret_last ? _GEN_828 : dirty_0_95; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1346 = ret_last ? _GEN_829 : dirty_0_96; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1347 = ret_last ? _GEN_830 : dirty_0_97; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1348 = ret_last ? _GEN_831 : dirty_0_98; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1349 = ret_last ? _GEN_832 : dirty_0_99; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1350 = ret_last ? _GEN_833 : dirty_0_100; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1351 = ret_last ? _GEN_834 : dirty_0_101; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1352 = ret_last ? _GEN_835 : dirty_0_102; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1353 = ret_last ? _GEN_836 : dirty_0_103; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1354 = ret_last ? _GEN_837 : dirty_0_104; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1355 = ret_last ? _GEN_838 : dirty_0_105; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1356 = ret_last ? _GEN_839 : dirty_0_106; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1357 = ret_last ? _GEN_840 : dirty_0_107; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1358 = ret_last ? _GEN_841 : dirty_0_108; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1359 = ret_last ? _GEN_842 : dirty_0_109; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1360 = ret_last ? _GEN_843 : dirty_0_110; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1361 = ret_last ? _GEN_844 : dirty_0_111; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1362 = ret_last ? _GEN_845 : dirty_0_112; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1363 = ret_last ? _GEN_846 : dirty_0_113; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1364 = ret_last ? _GEN_847 : dirty_0_114; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1365 = ret_last ? _GEN_848 : dirty_0_115; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1366 = ret_last ? _GEN_849 : dirty_0_116; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1367 = ret_last ? _GEN_850 : dirty_0_117; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1368 = ret_last ? _GEN_851 : dirty_0_118; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1369 = ret_last ? _GEN_852 : dirty_0_119; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1370 = ret_last ? _GEN_853 : dirty_0_120; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1371 = ret_last ? _GEN_854 : dirty_0_121; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1372 = ret_last ? _GEN_855 : dirty_0_122; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1373 = ret_last ? _GEN_856 : dirty_0_123; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1374 = ret_last ? _GEN_857 : dirty_0_124; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1375 = ret_last ? _GEN_858 : dirty_0_125; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1376 = ret_last ? _GEN_859 : dirty_0_126; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1377 = ret_last ? _GEN_860 : dirty_0_127; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1378 = ret_last ? _GEN_861 : dirty_0_128; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1379 = ret_last ? _GEN_862 : dirty_0_129; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1380 = ret_last ? _GEN_863 : dirty_0_130; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1381 = ret_last ? _GEN_864 : dirty_0_131; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1382 = ret_last ? _GEN_865 : dirty_0_132; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1383 = ret_last ? _GEN_866 : dirty_0_133; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1384 = ret_last ? _GEN_867 : dirty_0_134; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1385 = ret_last ? _GEN_868 : dirty_0_135; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1386 = ret_last ? _GEN_869 : dirty_0_136; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1387 = ret_last ? _GEN_870 : dirty_0_137; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1388 = ret_last ? _GEN_871 : dirty_0_138; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1389 = ret_last ? _GEN_872 : dirty_0_139; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1390 = ret_last ? _GEN_873 : dirty_0_140; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1391 = ret_last ? _GEN_874 : dirty_0_141; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1392 = ret_last ? _GEN_875 : dirty_0_142; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1393 = ret_last ? _GEN_876 : dirty_0_143; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1394 = ret_last ? _GEN_877 : dirty_0_144; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1395 = ret_last ? _GEN_878 : dirty_0_145; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1396 = ret_last ? _GEN_879 : dirty_0_146; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1397 = ret_last ? _GEN_880 : dirty_0_147; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1398 = ret_last ? _GEN_881 : dirty_0_148; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1399 = ret_last ? _GEN_882 : dirty_0_149; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1400 = ret_last ? _GEN_883 : dirty_0_150; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1401 = ret_last ? _GEN_884 : dirty_0_151; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1402 = ret_last ? _GEN_885 : dirty_0_152; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1403 = ret_last ? _GEN_886 : dirty_0_153; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1404 = ret_last ? _GEN_887 : dirty_0_154; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1405 = ret_last ? _GEN_888 : dirty_0_155; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1406 = ret_last ? _GEN_889 : dirty_0_156; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1407 = ret_last ? _GEN_890 : dirty_0_157; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1408 = ret_last ? _GEN_891 : dirty_0_158; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1409 = ret_last ? _GEN_892 : dirty_0_159; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1410 = ret_last ? _GEN_893 : dirty_0_160; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1411 = ret_last ? _GEN_894 : dirty_0_161; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1412 = ret_last ? _GEN_895 : dirty_0_162; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1413 = ret_last ? _GEN_896 : dirty_0_163; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1414 = ret_last ? _GEN_897 : dirty_0_164; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1415 = ret_last ? _GEN_898 : dirty_0_165; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1416 = ret_last ? _GEN_899 : dirty_0_166; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1417 = ret_last ? _GEN_900 : dirty_0_167; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1418 = ret_last ? _GEN_901 : dirty_0_168; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1419 = ret_last ? _GEN_902 : dirty_0_169; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1420 = ret_last ? _GEN_903 : dirty_0_170; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1421 = ret_last ? _GEN_904 : dirty_0_171; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1422 = ret_last ? _GEN_905 : dirty_0_172; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1423 = ret_last ? _GEN_906 : dirty_0_173; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1424 = ret_last ? _GEN_907 : dirty_0_174; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1425 = ret_last ? _GEN_908 : dirty_0_175; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1426 = ret_last ? _GEN_909 : dirty_0_176; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1427 = ret_last ? _GEN_910 : dirty_0_177; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1428 = ret_last ? _GEN_911 : dirty_0_178; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1429 = ret_last ? _GEN_912 : dirty_0_179; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1430 = ret_last ? _GEN_913 : dirty_0_180; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1431 = ret_last ? _GEN_914 : dirty_0_181; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1432 = ret_last ? _GEN_915 : dirty_0_182; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1433 = ret_last ? _GEN_916 : dirty_0_183; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1434 = ret_last ? _GEN_917 : dirty_0_184; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1435 = ret_last ? _GEN_918 : dirty_0_185; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1436 = ret_last ? _GEN_919 : dirty_0_186; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1437 = ret_last ? _GEN_920 : dirty_0_187; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1438 = ret_last ? _GEN_921 : dirty_0_188; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1439 = ret_last ? _GEN_922 : dirty_0_189; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1440 = ret_last ? _GEN_923 : dirty_0_190; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1441 = ret_last ? _GEN_924 : dirty_0_191; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1442 = ret_last ? _GEN_925 : dirty_0_192; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1443 = ret_last ? _GEN_926 : dirty_0_193; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1444 = ret_last ? _GEN_927 : dirty_0_194; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1445 = ret_last ? _GEN_928 : dirty_0_195; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1446 = ret_last ? _GEN_929 : dirty_0_196; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1447 = ret_last ? _GEN_930 : dirty_0_197; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1448 = ret_last ? _GEN_931 : dirty_0_198; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1449 = ret_last ? _GEN_932 : dirty_0_199; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1450 = ret_last ? _GEN_933 : dirty_0_200; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1451 = ret_last ? _GEN_934 : dirty_0_201; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1452 = ret_last ? _GEN_935 : dirty_0_202; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1453 = ret_last ? _GEN_936 : dirty_0_203; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1454 = ret_last ? _GEN_937 : dirty_0_204; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1455 = ret_last ? _GEN_938 : dirty_0_205; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1456 = ret_last ? _GEN_939 : dirty_0_206; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1457 = ret_last ? _GEN_940 : dirty_0_207; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1458 = ret_last ? _GEN_941 : dirty_0_208; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1459 = ret_last ? _GEN_942 : dirty_0_209; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1460 = ret_last ? _GEN_943 : dirty_0_210; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1461 = ret_last ? _GEN_944 : dirty_0_211; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1462 = ret_last ? _GEN_945 : dirty_0_212; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1463 = ret_last ? _GEN_946 : dirty_0_213; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1464 = ret_last ? _GEN_947 : dirty_0_214; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1465 = ret_last ? _GEN_948 : dirty_0_215; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1466 = ret_last ? _GEN_949 : dirty_0_216; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1467 = ret_last ? _GEN_950 : dirty_0_217; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1468 = ret_last ? _GEN_951 : dirty_0_218; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1469 = ret_last ? _GEN_952 : dirty_0_219; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1470 = ret_last ? _GEN_953 : dirty_0_220; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1471 = ret_last ? _GEN_954 : dirty_0_221; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1472 = ret_last ? _GEN_955 : dirty_0_222; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1473 = ret_last ? _GEN_956 : dirty_0_223; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1474 = ret_last ? _GEN_957 : dirty_0_224; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1475 = ret_last ? _GEN_958 : dirty_0_225; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1476 = ret_last ? _GEN_959 : dirty_0_226; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1477 = ret_last ? _GEN_960 : dirty_0_227; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1478 = ret_last ? _GEN_961 : dirty_0_228; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1479 = ret_last ? _GEN_962 : dirty_0_229; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1480 = ret_last ? _GEN_963 : dirty_0_230; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1481 = ret_last ? _GEN_964 : dirty_0_231; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1482 = ret_last ? _GEN_965 : dirty_0_232; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1483 = ret_last ? _GEN_966 : dirty_0_233; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1484 = ret_last ? _GEN_967 : dirty_0_234; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1485 = ret_last ? _GEN_968 : dirty_0_235; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1486 = ret_last ? _GEN_969 : dirty_0_236; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1487 = ret_last ? _GEN_970 : dirty_0_237; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1488 = ret_last ? _GEN_971 : dirty_0_238; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1489 = ret_last ? _GEN_972 : dirty_0_239; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1490 = ret_last ? _GEN_973 : dirty_0_240; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1491 = ret_last ? _GEN_974 : dirty_0_241; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1492 = ret_last ? _GEN_975 : dirty_0_242; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1493 = ret_last ? _GEN_976 : dirty_0_243; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1494 = ret_last ? _GEN_977 : dirty_0_244; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1495 = ret_last ? _GEN_978 : dirty_0_245; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1496 = ret_last ? _GEN_979 : dirty_0_246; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1497 = ret_last ? _GEN_980 : dirty_0_247; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1498 = ret_last ? _GEN_981 : dirty_0_248; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1499 = ret_last ? _GEN_982 : dirty_0_249; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1500 = ret_last ? _GEN_983 : dirty_0_250; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1501 = ret_last ? _GEN_984 : dirty_0_251; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1502 = ret_last ? _GEN_985 : dirty_0_252; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1503 = ret_last ? _GEN_986 : dirty_0_253; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1504 = ret_last ? _GEN_987 : dirty_0_254; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1505 = ret_last ? _GEN_988 : dirty_0_255; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1506 = ret_last ? _GEN_989 : dirty_1_0; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1507 = ret_last ? _GEN_990 : dirty_1_1; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1508 = ret_last ? _GEN_991 : dirty_1_2; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1509 = ret_last ? _GEN_992 : dirty_1_3; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1510 = ret_last ? _GEN_993 : dirty_1_4; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1511 = ret_last ? _GEN_994 : dirty_1_5; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1512 = ret_last ? _GEN_995 : dirty_1_6; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1513 = ret_last ? _GEN_996 : dirty_1_7; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1514 = ret_last ? _GEN_997 : dirty_1_8; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1515 = ret_last ? _GEN_998 : dirty_1_9; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1516 = ret_last ? _GEN_999 : dirty_1_10; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1517 = ret_last ? _GEN_1000 : dirty_1_11; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1518 = ret_last ? _GEN_1001 : dirty_1_12; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1519 = ret_last ? _GEN_1002 : dirty_1_13; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1520 = ret_last ? _GEN_1003 : dirty_1_14; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1521 = ret_last ? _GEN_1004 : dirty_1_15; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1522 = ret_last ? _GEN_1005 : dirty_1_16; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1523 = ret_last ? _GEN_1006 : dirty_1_17; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1524 = ret_last ? _GEN_1007 : dirty_1_18; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1525 = ret_last ? _GEN_1008 : dirty_1_19; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1526 = ret_last ? _GEN_1009 : dirty_1_20; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1527 = ret_last ? _GEN_1010 : dirty_1_21; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1528 = ret_last ? _GEN_1011 : dirty_1_22; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1529 = ret_last ? _GEN_1012 : dirty_1_23; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1530 = ret_last ? _GEN_1013 : dirty_1_24; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1531 = ret_last ? _GEN_1014 : dirty_1_25; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1532 = ret_last ? _GEN_1015 : dirty_1_26; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1533 = ret_last ? _GEN_1016 : dirty_1_27; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1534 = ret_last ? _GEN_1017 : dirty_1_28; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1535 = ret_last ? _GEN_1018 : dirty_1_29; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1536 = ret_last ? _GEN_1019 : dirty_1_30; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1537 = ret_last ? _GEN_1020 : dirty_1_31; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1538 = ret_last ? _GEN_1021 : dirty_1_32; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1539 = ret_last ? _GEN_1022 : dirty_1_33; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1540 = ret_last ? _GEN_1023 : dirty_1_34; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1541 = ret_last ? _GEN_1024 : dirty_1_35; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1542 = ret_last ? _GEN_1025 : dirty_1_36; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1543 = ret_last ? _GEN_1026 : dirty_1_37; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1544 = ret_last ? _GEN_1027 : dirty_1_38; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1545 = ret_last ? _GEN_1028 : dirty_1_39; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1546 = ret_last ? _GEN_1029 : dirty_1_40; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1547 = ret_last ? _GEN_1030 : dirty_1_41; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1548 = ret_last ? _GEN_1031 : dirty_1_42; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1549 = ret_last ? _GEN_1032 : dirty_1_43; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1550 = ret_last ? _GEN_1033 : dirty_1_44; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1551 = ret_last ? _GEN_1034 : dirty_1_45; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1552 = ret_last ? _GEN_1035 : dirty_1_46; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1553 = ret_last ? _GEN_1036 : dirty_1_47; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1554 = ret_last ? _GEN_1037 : dirty_1_48; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1555 = ret_last ? _GEN_1038 : dirty_1_49; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1556 = ret_last ? _GEN_1039 : dirty_1_50; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1557 = ret_last ? _GEN_1040 : dirty_1_51; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1558 = ret_last ? _GEN_1041 : dirty_1_52; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1559 = ret_last ? _GEN_1042 : dirty_1_53; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1560 = ret_last ? _GEN_1043 : dirty_1_54; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1561 = ret_last ? _GEN_1044 : dirty_1_55; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1562 = ret_last ? _GEN_1045 : dirty_1_56; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1563 = ret_last ? _GEN_1046 : dirty_1_57; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1564 = ret_last ? _GEN_1047 : dirty_1_58; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1565 = ret_last ? _GEN_1048 : dirty_1_59; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1566 = ret_last ? _GEN_1049 : dirty_1_60; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1567 = ret_last ? _GEN_1050 : dirty_1_61; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1568 = ret_last ? _GEN_1051 : dirty_1_62; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1569 = ret_last ? _GEN_1052 : dirty_1_63; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1570 = ret_last ? _GEN_1053 : dirty_1_64; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1571 = ret_last ? _GEN_1054 : dirty_1_65; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1572 = ret_last ? _GEN_1055 : dirty_1_66; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1573 = ret_last ? _GEN_1056 : dirty_1_67; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1574 = ret_last ? _GEN_1057 : dirty_1_68; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1575 = ret_last ? _GEN_1058 : dirty_1_69; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1576 = ret_last ? _GEN_1059 : dirty_1_70; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1577 = ret_last ? _GEN_1060 : dirty_1_71; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1578 = ret_last ? _GEN_1061 : dirty_1_72; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1579 = ret_last ? _GEN_1062 : dirty_1_73; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1580 = ret_last ? _GEN_1063 : dirty_1_74; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1581 = ret_last ? _GEN_1064 : dirty_1_75; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1582 = ret_last ? _GEN_1065 : dirty_1_76; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1583 = ret_last ? _GEN_1066 : dirty_1_77; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1584 = ret_last ? _GEN_1067 : dirty_1_78; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1585 = ret_last ? _GEN_1068 : dirty_1_79; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1586 = ret_last ? _GEN_1069 : dirty_1_80; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1587 = ret_last ? _GEN_1070 : dirty_1_81; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1588 = ret_last ? _GEN_1071 : dirty_1_82; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1589 = ret_last ? _GEN_1072 : dirty_1_83; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1590 = ret_last ? _GEN_1073 : dirty_1_84; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1591 = ret_last ? _GEN_1074 : dirty_1_85; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1592 = ret_last ? _GEN_1075 : dirty_1_86; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1593 = ret_last ? _GEN_1076 : dirty_1_87; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1594 = ret_last ? _GEN_1077 : dirty_1_88; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1595 = ret_last ? _GEN_1078 : dirty_1_89; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1596 = ret_last ? _GEN_1079 : dirty_1_90; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1597 = ret_last ? _GEN_1080 : dirty_1_91; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1598 = ret_last ? _GEN_1081 : dirty_1_92; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1599 = ret_last ? _GEN_1082 : dirty_1_93; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1600 = ret_last ? _GEN_1083 : dirty_1_94; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1601 = ret_last ? _GEN_1084 : dirty_1_95; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1602 = ret_last ? _GEN_1085 : dirty_1_96; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1603 = ret_last ? _GEN_1086 : dirty_1_97; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1604 = ret_last ? _GEN_1087 : dirty_1_98; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1605 = ret_last ? _GEN_1088 : dirty_1_99; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1606 = ret_last ? _GEN_1089 : dirty_1_100; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1607 = ret_last ? _GEN_1090 : dirty_1_101; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1608 = ret_last ? _GEN_1091 : dirty_1_102; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1609 = ret_last ? _GEN_1092 : dirty_1_103; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1610 = ret_last ? _GEN_1093 : dirty_1_104; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1611 = ret_last ? _GEN_1094 : dirty_1_105; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1612 = ret_last ? _GEN_1095 : dirty_1_106; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1613 = ret_last ? _GEN_1096 : dirty_1_107; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1614 = ret_last ? _GEN_1097 : dirty_1_108; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1615 = ret_last ? _GEN_1098 : dirty_1_109; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1616 = ret_last ? _GEN_1099 : dirty_1_110; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1617 = ret_last ? _GEN_1100 : dirty_1_111; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1618 = ret_last ? _GEN_1101 : dirty_1_112; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1619 = ret_last ? _GEN_1102 : dirty_1_113; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1620 = ret_last ? _GEN_1103 : dirty_1_114; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1621 = ret_last ? _GEN_1104 : dirty_1_115; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1622 = ret_last ? _GEN_1105 : dirty_1_116; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1623 = ret_last ? _GEN_1106 : dirty_1_117; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1624 = ret_last ? _GEN_1107 : dirty_1_118; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1625 = ret_last ? _GEN_1108 : dirty_1_119; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1626 = ret_last ? _GEN_1109 : dirty_1_120; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1627 = ret_last ? _GEN_1110 : dirty_1_121; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1628 = ret_last ? _GEN_1111 : dirty_1_122; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1629 = ret_last ? _GEN_1112 : dirty_1_123; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1630 = ret_last ? _GEN_1113 : dirty_1_124; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1631 = ret_last ? _GEN_1114 : dirty_1_125; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1632 = ret_last ? _GEN_1115 : dirty_1_126; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1633 = ret_last ? _GEN_1116 : dirty_1_127; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1634 = ret_last ? _GEN_1117 : dirty_1_128; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1635 = ret_last ? _GEN_1118 : dirty_1_129; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1636 = ret_last ? _GEN_1119 : dirty_1_130; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1637 = ret_last ? _GEN_1120 : dirty_1_131; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1638 = ret_last ? _GEN_1121 : dirty_1_132; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1639 = ret_last ? _GEN_1122 : dirty_1_133; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1640 = ret_last ? _GEN_1123 : dirty_1_134; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1641 = ret_last ? _GEN_1124 : dirty_1_135; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1642 = ret_last ? _GEN_1125 : dirty_1_136; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1643 = ret_last ? _GEN_1126 : dirty_1_137; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1644 = ret_last ? _GEN_1127 : dirty_1_138; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1645 = ret_last ? _GEN_1128 : dirty_1_139; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1646 = ret_last ? _GEN_1129 : dirty_1_140; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1647 = ret_last ? _GEN_1130 : dirty_1_141; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1648 = ret_last ? _GEN_1131 : dirty_1_142; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1649 = ret_last ? _GEN_1132 : dirty_1_143; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1650 = ret_last ? _GEN_1133 : dirty_1_144; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1651 = ret_last ? _GEN_1134 : dirty_1_145; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1652 = ret_last ? _GEN_1135 : dirty_1_146; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1653 = ret_last ? _GEN_1136 : dirty_1_147; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1654 = ret_last ? _GEN_1137 : dirty_1_148; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1655 = ret_last ? _GEN_1138 : dirty_1_149; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1656 = ret_last ? _GEN_1139 : dirty_1_150; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1657 = ret_last ? _GEN_1140 : dirty_1_151; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1658 = ret_last ? _GEN_1141 : dirty_1_152; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1659 = ret_last ? _GEN_1142 : dirty_1_153; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1660 = ret_last ? _GEN_1143 : dirty_1_154; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1661 = ret_last ? _GEN_1144 : dirty_1_155; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1662 = ret_last ? _GEN_1145 : dirty_1_156; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1663 = ret_last ? _GEN_1146 : dirty_1_157; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1664 = ret_last ? _GEN_1147 : dirty_1_158; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1665 = ret_last ? _GEN_1148 : dirty_1_159; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1666 = ret_last ? _GEN_1149 : dirty_1_160; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1667 = ret_last ? _GEN_1150 : dirty_1_161; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1668 = ret_last ? _GEN_1151 : dirty_1_162; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1669 = ret_last ? _GEN_1152 : dirty_1_163; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1670 = ret_last ? _GEN_1153 : dirty_1_164; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1671 = ret_last ? _GEN_1154 : dirty_1_165; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1672 = ret_last ? _GEN_1155 : dirty_1_166; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1673 = ret_last ? _GEN_1156 : dirty_1_167; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1674 = ret_last ? _GEN_1157 : dirty_1_168; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1675 = ret_last ? _GEN_1158 : dirty_1_169; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1676 = ret_last ? _GEN_1159 : dirty_1_170; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1677 = ret_last ? _GEN_1160 : dirty_1_171; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1678 = ret_last ? _GEN_1161 : dirty_1_172; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1679 = ret_last ? _GEN_1162 : dirty_1_173; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1680 = ret_last ? _GEN_1163 : dirty_1_174; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1681 = ret_last ? _GEN_1164 : dirty_1_175; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1682 = ret_last ? _GEN_1165 : dirty_1_176; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1683 = ret_last ? _GEN_1166 : dirty_1_177; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1684 = ret_last ? _GEN_1167 : dirty_1_178; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1685 = ret_last ? _GEN_1168 : dirty_1_179; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1686 = ret_last ? _GEN_1169 : dirty_1_180; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1687 = ret_last ? _GEN_1170 : dirty_1_181; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1688 = ret_last ? _GEN_1171 : dirty_1_182; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1689 = ret_last ? _GEN_1172 : dirty_1_183; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1690 = ret_last ? _GEN_1173 : dirty_1_184; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1691 = ret_last ? _GEN_1174 : dirty_1_185; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1692 = ret_last ? _GEN_1175 : dirty_1_186; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1693 = ret_last ? _GEN_1176 : dirty_1_187; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1694 = ret_last ? _GEN_1177 : dirty_1_188; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1695 = ret_last ? _GEN_1178 : dirty_1_189; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1696 = ret_last ? _GEN_1179 : dirty_1_190; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1697 = ret_last ? _GEN_1180 : dirty_1_191; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1698 = ret_last ? _GEN_1181 : dirty_1_192; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1699 = ret_last ? _GEN_1182 : dirty_1_193; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1700 = ret_last ? _GEN_1183 : dirty_1_194; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1701 = ret_last ? _GEN_1184 : dirty_1_195; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1702 = ret_last ? _GEN_1185 : dirty_1_196; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1703 = ret_last ? _GEN_1186 : dirty_1_197; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1704 = ret_last ? _GEN_1187 : dirty_1_198; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1705 = ret_last ? _GEN_1188 : dirty_1_199; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1706 = ret_last ? _GEN_1189 : dirty_1_200; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1707 = ret_last ? _GEN_1190 : dirty_1_201; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1708 = ret_last ? _GEN_1191 : dirty_1_202; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1709 = ret_last ? _GEN_1192 : dirty_1_203; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1710 = ret_last ? _GEN_1193 : dirty_1_204; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1711 = ret_last ? _GEN_1194 : dirty_1_205; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1712 = ret_last ? _GEN_1195 : dirty_1_206; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1713 = ret_last ? _GEN_1196 : dirty_1_207; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1714 = ret_last ? _GEN_1197 : dirty_1_208; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1715 = ret_last ? _GEN_1198 : dirty_1_209; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1716 = ret_last ? _GEN_1199 : dirty_1_210; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1717 = ret_last ? _GEN_1200 : dirty_1_211; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1718 = ret_last ? _GEN_1201 : dirty_1_212; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1719 = ret_last ? _GEN_1202 : dirty_1_213; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1720 = ret_last ? _GEN_1203 : dirty_1_214; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1721 = ret_last ? _GEN_1204 : dirty_1_215; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1722 = ret_last ? _GEN_1205 : dirty_1_216; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1723 = ret_last ? _GEN_1206 : dirty_1_217; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1724 = ret_last ? _GEN_1207 : dirty_1_218; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1725 = ret_last ? _GEN_1208 : dirty_1_219; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1726 = ret_last ? _GEN_1209 : dirty_1_220; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1727 = ret_last ? _GEN_1210 : dirty_1_221; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1728 = ret_last ? _GEN_1211 : dirty_1_222; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1729 = ret_last ? _GEN_1212 : dirty_1_223; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1730 = ret_last ? _GEN_1213 : dirty_1_224; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1731 = ret_last ? _GEN_1214 : dirty_1_225; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1732 = ret_last ? _GEN_1215 : dirty_1_226; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1733 = ret_last ? _GEN_1216 : dirty_1_227; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1734 = ret_last ? _GEN_1217 : dirty_1_228; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1735 = ret_last ? _GEN_1218 : dirty_1_229; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1736 = ret_last ? _GEN_1219 : dirty_1_230; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1737 = ret_last ? _GEN_1220 : dirty_1_231; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1738 = ret_last ? _GEN_1221 : dirty_1_232; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1739 = ret_last ? _GEN_1222 : dirty_1_233; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1740 = ret_last ? _GEN_1223 : dirty_1_234; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1741 = ret_last ? _GEN_1224 : dirty_1_235; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1742 = ret_last ? _GEN_1225 : dirty_1_236; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1743 = ret_last ? _GEN_1226 : dirty_1_237; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1744 = ret_last ? _GEN_1227 : dirty_1_238; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1745 = ret_last ? _GEN_1228 : dirty_1_239; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1746 = ret_last ? _GEN_1229 : dirty_1_240; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1747 = ret_last ? _GEN_1230 : dirty_1_241; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1748 = ret_last ? _GEN_1231 : dirty_1_242; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1749 = ret_last ? _GEN_1232 : dirty_1_243; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1750 = ret_last ? _GEN_1233 : dirty_1_244; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1751 = ret_last ? _GEN_1234 : dirty_1_245; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1752 = ret_last ? _GEN_1235 : dirty_1_246; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1753 = ret_last ? _GEN_1236 : dirty_1_247; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1754 = ret_last ? _GEN_1237 : dirty_1_248; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1755 = ret_last ? _GEN_1238 : dirty_1_249; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1756 = ret_last ? _GEN_1239 : dirty_1_250; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1757 = ret_last ? _GEN_1240 : dirty_1_251; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1758 = ret_last ? _GEN_1241 : dirty_1_252; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1759 = ret_last ? _GEN_1242 : dirty_1_253; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1760 = ret_last ? _GEN_1243 : dirty_1_254; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1761 = ret_last ? _GEN_1244 : dirty_1_255; // @[dcache.scala 389:21 113:28]
  wire  _GEN_1762 = ret_last & _GEN_11958; // @[dcache.scala 389:21 144:25]
  wire  _GEN_1763 = ret_last & refillIDX_r; // @[dcache.scala 389:21 144:25]
  wire [20:0] _GEN_1764 = ret_last ? _GEN_1247 : 21'h0; // @[dcache.scala 389:21 143:25]
  wire [20:0] _GEN_1765 = ret_last ? _GEN_1248 : 21'h0; // @[dcache.scala 389:21 143:25]
  wire [1:0] _GEN_1766 = ret_valid ? _wr_cnt_T_1 : wr_cnt; // @[dcache.scala 384:17 178:34 385:61]
  wire [31:0] _GEN_1767 = ret_valid ? _GEN_717 : 32'h0; // @[dcache.scala 384:17 149:33]
  wire [31:0] _GEN_1768 = ret_valid ? _GEN_718 : 32'h0; // @[dcache.scala 384:17 149:33]
  wire [31:0] _GEN_1769 = ret_valid ? _GEN_719 : 32'h0; // @[dcache.scala 384:17 149:33]
  wire [31:0] _GEN_1770 = ret_valid ? _GEN_720 : 32'h0; // @[dcache.scala 384:17 149:33]
  wire [31:0] _GEN_1771 = ret_valid ? _GEN_721 : 32'h0; // @[dcache.scala 384:17 149:33]
  wire [31:0] _GEN_1772 = ret_valid ? _GEN_722 : 32'h0; // @[dcache.scala 384:17 149:33]
  wire [31:0] _GEN_1773 = ret_valid ? _GEN_723 : 32'h0; // @[dcache.scala 384:17 149:33]
  wire [31:0] _GEN_1774 = ret_valid ? _GEN_724 : 32'h0; // @[dcache.scala 384:17 149:33]
  wire [3:0] _GEN_1775 = ret_valid ? _GEN_725 : 4'h0; // @[dcache.scala 384:17 150:33]
  wire [3:0] _GEN_1776 = ret_valid ? _GEN_726 : 4'h0; // @[dcache.scala 384:17 150:33]
  wire [3:0] _GEN_1777 = ret_valid ? _GEN_727 : 4'h0; // @[dcache.scala 384:17 150:33]
  wire [3:0] _GEN_1778 = ret_valid ? _GEN_728 : 4'h0; // @[dcache.scala 384:17 150:33]
  wire [3:0] _GEN_1779 = ret_valid ? _GEN_729 : 4'h0; // @[dcache.scala 384:17 150:33]
  wire [3:0] _GEN_1780 = ret_valid ? _GEN_730 : 4'h0; // @[dcache.scala 384:17 150:33]
  wire [3:0] _GEN_1781 = ret_valid ? _GEN_731 : 4'h0; // @[dcache.scala 384:17 150:33]
  wire [3:0] _GEN_1782 = ret_valid ? _GEN_732 : 4'h0; // @[dcache.scala 384:17 150:33]
  wire [2:0] _GEN_1783 = ret_valid ? _GEN_1249 : 3'h5; // @[dcache.scala 384:17 380:41]
  wire  _GEN_1784 = ret_valid ? _GEN_1250 : dirty_0_0; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1785 = ret_valid ? _GEN_1251 : dirty_0_1; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1786 = ret_valid ? _GEN_1252 : dirty_0_2; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1787 = ret_valid ? _GEN_1253 : dirty_0_3; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1788 = ret_valid ? _GEN_1254 : dirty_0_4; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1789 = ret_valid ? _GEN_1255 : dirty_0_5; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1790 = ret_valid ? _GEN_1256 : dirty_0_6; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1791 = ret_valid ? _GEN_1257 : dirty_0_7; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1792 = ret_valid ? _GEN_1258 : dirty_0_8; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1793 = ret_valid ? _GEN_1259 : dirty_0_9; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1794 = ret_valid ? _GEN_1260 : dirty_0_10; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1795 = ret_valid ? _GEN_1261 : dirty_0_11; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1796 = ret_valid ? _GEN_1262 : dirty_0_12; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1797 = ret_valid ? _GEN_1263 : dirty_0_13; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1798 = ret_valid ? _GEN_1264 : dirty_0_14; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1799 = ret_valid ? _GEN_1265 : dirty_0_15; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1800 = ret_valid ? _GEN_1266 : dirty_0_16; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1801 = ret_valid ? _GEN_1267 : dirty_0_17; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1802 = ret_valid ? _GEN_1268 : dirty_0_18; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1803 = ret_valid ? _GEN_1269 : dirty_0_19; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1804 = ret_valid ? _GEN_1270 : dirty_0_20; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1805 = ret_valid ? _GEN_1271 : dirty_0_21; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1806 = ret_valid ? _GEN_1272 : dirty_0_22; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1807 = ret_valid ? _GEN_1273 : dirty_0_23; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1808 = ret_valid ? _GEN_1274 : dirty_0_24; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1809 = ret_valid ? _GEN_1275 : dirty_0_25; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1810 = ret_valid ? _GEN_1276 : dirty_0_26; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1811 = ret_valid ? _GEN_1277 : dirty_0_27; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1812 = ret_valid ? _GEN_1278 : dirty_0_28; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1813 = ret_valid ? _GEN_1279 : dirty_0_29; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1814 = ret_valid ? _GEN_1280 : dirty_0_30; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1815 = ret_valid ? _GEN_1281 : dirty_0_31; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1816 = ret_valid ? _GEN_1282 : dirty_0_32; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1817 = ret_valid ? _GEN_1283 : dirty_0_33; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1818 = ret_valid ? _GEN_1284 : dirty_0_34; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1819 = ret_valid ? _GEN_1285 : dirty_0_35; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1820 = ret_valid ? _GEN_1286 : dirty_0_36; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1821 = ret_valid ? _GEN_1287 : dirty_0_37; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1822 = ret_valid ? _GEN_1288 : dirty_0_38; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1823 = ret_valid ? _GEN_1289 : dirty_0_39; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1824 = ret_valid ? _GEN_1290 : dirty_0_40; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1825 = ret_valid ? _GEN_1291 : dirty_0_41; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1826 = ret_valid ? _GEN_1292 : dirty_0_42; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1827 = ret_valid ? _GEN_1293 : dirty_0_43; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1828 = ret_valid ? _GEN_1294 : dirty_0_44; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1829 = ret_valid ? _GEN_1295 : dirty_0_45; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1830 = ret_valid ? _GEN_1296 : dirty_0_46; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1831 = ret_valid ? _GEN_1297 : dirty_0_47; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1832 = ret_valid ? _GEN_1298 : dirty_0_48; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1833 = ret_valid ? _GEN_1299 : dirty_0_49; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1834 = ret_valid ? _GEN_1300 : dirty_0_50; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1835 = ret_valid ? _GEN_1301 : dirty_0_51; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1836 = ret_valid ? _GEN_1302 : dirty_0_52; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1837 = ret_valid ? _GEN_1303 : dirty_0_53; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1838 = ret_valid ? _GEN_1304 : dirty_0_54; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1839 = ret_valid ? _GEN_1305 : dirty_0_55; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1840 = ret_valid ? _GEN_1306 : dirty_0_56; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1841 = ret_valid ? _GEN_1307 : dirty_0_57; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1842 = ret_valid ? _GEN_1308 : dirty_0_58; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1843 = ret_valid ? _GEN_1309 : dirty_0_59; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1844 = ret_valid ? _GEN_1310 : dirty_0_60; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1845 = ret_valid ? _GEN_1311 : dirty_0_61; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1846 = ret_valid ? _GEN_1312 : dirty_0_62; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1847 = ret_valid ? _GEN_1313 : dirty_0_63; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1848 = ret_valid ? _GEN_1314 : dirty_0_64; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1849 = ret_valid ? _GEN_1315 : dirty_0_65; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1850 = ret_valid ? _GEN_1316 : dirty_0_66; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1851 = ret_valid ? _GEN_1317 : dirty_0_67; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1852 = ret_valid ? _GEN_1318 : dirty_0_68; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1853 = ret_valid ? _GEN_1319 : dirty_0_69; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1854 = ret_valid ? _GEN_1320 : dirty_0_70; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1855 = ret_valid ? _GEN_1321 : dirty_0_71; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1856 = ret_valid ? _GEN_1322 : dirty_0_72; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1857 = ret_valid ? _GEN_1323 : dirty_0_73; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1858 = ret_valid ? _GEN_1324 : dirty_0_74; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1859 = ret_valid ? _GEN_1325 : dirty_0_75; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1860 = ret_valid ? _GEN_1326 : dirty_0_76; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1861 = ret_valid ? _GEN_1327 : dirty_0_77; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1862 = ret_valid ? _GEN_1328 : dirty_0_78; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1863 = ret_valid ? _GEN_1329 : dirty_0_79; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1864 = ret_valid ? _GEN_1330 : dirty_0_80; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1865 = ret_valid ? _GEN_1331 : dirty_0_81; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1866 = ret_valid ? _GEN_1332 : dirty_0_82; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1867 = ret_valid ? _GEN_1333 : dirty_0_83; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1868 = ret_valid ? _GEN_1334 : dirty_0_84; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1869 = ret_valid ? _GEN_1335 : dirty_0_85; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1870 = ret_valid ? _GEN_1336 : dirty_0_86; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1871 = ret_valid ? _GEN_1337 : dirty_0_87; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1872 = ret_valid ? _GEN_1338 : dirty_0_88; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1873 = ret_valid ? _GEN_1339 : dirty_0_89; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1874 = ret_valid ? _GEN_1340 : dirty_0_90; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1875 = ret_valid ? _GEN_1341 : dirty_0_91; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1876 = ret_valid ? _GEN_1342 : dirty_0_92; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1877 = ret_valid ? _GEN_1343 : dirty_0_93; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1878 = ret_valid ? _GEN_1344 : dirty_0_94; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1879 = ret_valid ? _GEN_1345 : dirty_0_95; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1880 = ret_valid ? _GEN_1346 : dirty_0_96; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1881 = ret_valid ? _GEN_1347 : dirty_0_97; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1882 = ret_valid ? _GEN_1348 : dirty_0_98; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1883 = ret_valid ? _GEN_1349 : dirty_0_99; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1884 = ret_valid ? _GEN_1350 : dirty_0_100; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1885 = ret_valid ? _GEN_1351 : dirty_0_101; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1886 = ret_valid ? _GEN_1352 : dirty_0_102; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1887 = ret_valid ? _GEN_1353 : dirty_0_103; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1888 = ret_valid ? _GEN_1354 : dirty_0_104; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1889 = ret_valid ? _GEN_1355 : dirty_0_105; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1890 = ret_valid ? _GEN_1356 : dirty_0_106; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1891 = ret_valid ? _GEN_1357 : dirty_0_107; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1892 = ret_valid ? _GEN_1358 : dirty_0_108; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1893 = ret_valid ? _GEN_1359 : dirty_0_109; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1894 = ret_valid ? _GEN_1360 : dirty_0_110; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1895 = ret_valid ? _GEN_1361 : dirty_0_111; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1896 = ret_valid ? _GEN_1362 : dirty_0_112; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1897 = ret_valid ? _GEN_1363 : dirty_0_113; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1898 = ret_valid ? _GEN_1364 : dirty_0_114; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1899 = ret_valid ? _GEN_1365 : dirty_0_115; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1900 = ret_valid ? _GEN_1366 : dirty_0_116; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1901 = ret_valid ? _GEN_1367 : dirty_0_117; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1902 = ret_valid ? _GEN_1368 : dirty_0_118; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1903 = ret_valid ? _GEN_1369 : dirty_0_119; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1904 = ret_valid ? _GEN_1370 : dirty_0_120; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1905 = ret_valid ? _GEN_1371 : dirty_0_121; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1906 = ret_valid ? _GEN_1372 : dirty_0_122; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1907 = ret_valid ? _GEN_1373 : dirty_0_123; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1908 = ret_valid ? _GEN_1374 : dirty_0_124; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1909 = ret_valid ? _GEN_1375 : dirty_0_125; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1910 = ret_valid ? _GEN_1376 : dirty_0_126; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1911 = ret_valid ? _GEN_1377 : dirty_0_127; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1912 = ret_valid ? _GEN_1378 : dirty_0_128; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1913 = ret_valid ? _GEN_1379 : dirty_0_129; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1914 = ret_valid ? _GEN_1380 : dirty_0_130; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1915 = ret_valid ? _GEN_1381 : dirty_0_131; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1916 = ret_valid ? _GEN_1382 : dirty_0_132; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1917 = ret_valid ? _GEN_1383 : dirty_0_133; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1918 = ret_valid ? _GEN_1384 : dirty_0_134; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1919 = ret_valid ? _GEN_1385 : dirty_0_135; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1920 = ret_valid ? _GEN_1386 : dirty_0_136; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1921 = ret_valid ? _GEN_1387 : dirty_0_137; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1922 = ret_valid ? _GEN_1388 : dirty_0_138; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1923 = ret_valid ? _GEN_1389 : dirty_0_139; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1924 = ret_valid ? _GEN_1390 : dirty_0_140; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1925 = ret_valid ? _GEN_1391 : dirty_0_141; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1926 = ret_valid ? _GEN_1392 : dirty_0_142; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1927 = ret_valid ? _GEN_1393 : dirty_0_143; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1928 = ret_valid ? _GEN_1394 : dirty_0_144; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1929 = ret_valid ? _GEN_1395 : dirty_0_145; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1930 = ret_valid ? _GEN_1396 : dirty_0_146; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1931 = ret_valid ? _GEN_1397 : dirty_0_147; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1932 = ret_valid ? _GEN_1398 : dirty_0_148; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1933 = ret_valid ? _GEN_1399 : dirty_0_149; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1934 = ret_valid ? _GEN_1400 : dirty_0_150; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1935 = ret_valid ? _GEN_1401 : dirty_0_151; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1936 = ret_valid ? _GEN_1402 : dirty_0_152; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1937 = ret_valid ? _GEN_1403 : dirty_0_153; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1938 = ret_valid ? _GEN_1404 : dirty_0_154; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1939 = ret_valid ? _GEN_1405 : dirty_0_155; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1940 = ret_valid ? _GEN_1406 : dirty_0_156; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1941 = ret_valid ? _GEN_1407 : dirty_0_157; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1942 = ret_valid ? _GEN_1408 : dirty_0_158; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1943 = ret_valid ? _GEN_1409 : dirty_0_159; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1944 = ret_valid ? _GEN_1410 : dirty_0_160; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1945 = ret_valid ? _GEN_1411 : dirty_0_161; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1946 = ret_valid ? _GEN_1412 : dirty_0_162; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1947 = ret_valid ? _GEN_1413 : dirty_0_163; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1948 = ret_valid ? _GEN_1414 : dirty_0_164; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1949 = ret_valid ? _GEN_1415 : dirty_0_165; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1950 = ret_valid ? _GEN_1416 : dirty_0_166; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1951 = ret_valid ? _GEN_1417 : dirty_0_167; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1952 = ret_valid ? _GEN_1418 : dirty_0_168; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1953 = ret_valid ? _GEN_1419 : dirty_0_169; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1954 = ret_valid ? _GEN_1420 : dirty_0_170; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1955 = ret_valid ? _GEN_1421 : dirty_0_171; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1956 = ret_valid ? _GEN_1422 : dirty_0_172; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1957 = ret_valid ? _GEN_1423 : dirty_0_173; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1958 = ret_valid ? _GEN_1424 : dirty_0_174; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1959 = ret_valid ? _GEN_1425 : dirty_0_175; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1960 = ret_valid ? _GEN_1426 : dirty_0_176; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1961 = ret_valid ? _GEN_1427 : dirty_0_177; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1962 = ret_valid ? _GEN_1428 : dirty_0_178; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1963 = ret_valid ? _GEN_1429 : dirty_0_179; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1964 = ret_valid ? _GEN_1430 : dirty_0_180; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1965 = ret_valid ? _GEN_1431 : dirty_0_181; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1966 = ret_valid ? _GEN_1432 : dirty_0_182; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1967 = ret_valid ? _GEN_1433 : dirty_0_183; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1968 = ret_valid ? _GEN_1434 : dirty_0_184; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1969 = ret_valid ? _GEN_1435 : dirty_0_185; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1970 = ret_valid ? _GEN_1436 : dirty_0_186; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1971 = ret_valid ? _GEN_1437 : dirty_0_187; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1972 = ret_valid ? _GEN_1438 : dirty_0_188; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1973 = ret_valid ? _GEN_1439 : dirty_0_189; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1974 = ret_valid ? _GEN_1440 : dirty_0_190; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1975 = ret_valid ? _GEN_1441 : dirty_0_191; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1976 = ret_valid ? _GEN_1442 : dirty_0_192; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1977 = ret_valid ? _GEN_1443 : dirty_0_193; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1978 = ret_valid ? _GEN_1444 : dirty_0_194; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1979 = ret_valid ? _GEN_1445 : dirty_0_195; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1980 = ret_valid ? _GEN_1446 : dirty_0_196; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1981 = ret_valid ? _GEN_1447 : dirty_0_197; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1982 = ret_valid ? _GEN_1448 : dirty_0_198; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1983 = ret_valid ? _GEN_1449 : dirty_0_199; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1984 = ret_valid ? _GEN_1450 : dirty_0_200; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1985 = ret_valid ? _GEN_1451 : dirty_0_201; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1986 = ret_valid ? _GEN_1452 : dirty_0_202; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1987 = ret_valid ? _GEN_1453 : dirty_0_203; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1988 = ret_valid ? _GEN_1454 : dirty_0_204; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1989 = ret_valid ? _GEN_1455 : dirty_0_205; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1990 = ret_valid ? _GEN_1456 : dirty_0_206; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1991 = ret_valid ? _GEN_1457 : dirty_0_207; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1992 = ret_valid ? _GEN_1458 : dirty_0_208; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1993 = ret_valid ? _GEN_1459 : dirty_0_209; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1994 = ret_valid ? _GEN_1460 : dirty_0_210; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1995 = ret_valid ? _GEN_1461 : dirty_0_211; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1996 = ret_valid ? _GEN_1462 : dirty_0_212; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1997 = ret_valid ? _GEN_1463 : dirty_0_213; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1998 = ret_valid ? _GEN_1464 : dirty_0_214; // @[dcache.scala 384:17 113:28]
  wire  _GEN_1999 = ret_valid ? _GEN_1465 : dirty_0_215; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2000 = ret_valid ? _GEN_1466 : dirty_0_216; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2001 = ret_valid ? _GEN_1467 : dirty_0_217; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2002 = ret_valid ? _GEN_1468 : dirty_0_218; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2003 = ret_valid ? _GEN_1469 : dirty_0_219; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2004 = ret_valid ? _GEN_1470 : dirty_0_220; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2005 = ret_valid ? _GEN_1471 : dirty_0_221; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2006 = ret_valid ? _GEN_1472 : dirty_0_222; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2007 = ret_valid ? _GEN_1473 : dirty_0_223; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2008 = ret_valid ? _GEN_1474 : dirty_0_224; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2009 = ret_valid ? _GEN_1475 : dirty_0_225; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2010 = ret_valid ? _GEN_1476 : dirty_0_226; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2011 = ret_valid ? _GEN_1477 : dirty_0_227; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2012 = ret_valid ? _GEN_1478 : dirty_0_228; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2013 = ret_valid ? _GEN_1479 : dirty_0_229; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2014 = ret_valid ? _GEN_1480 : dirty_0_230; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2015 = ret_valid ? _GEN_1481 : dirty_0_231; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2016 = ret_valid ? _GEN_1482 : dirty_0_232; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2017 = ret_valid ? _GEN_1483 : dirty_0_233; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2018 = ret_valid ? _GEN_1484 : dirty_0_234; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2019 = ret_valid ? _GEN_1485 : dirty_0_235; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2020 = ret_valid ? _GEN_1486 : dirty_0_236; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2021 = ret_valid ? _GEN_1487 : dirty_0_237; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2022 = ret_valid ? _GEN_1488 : dirty_0_238; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2023 = ret_valid ? _GEN_1489 : dirty_0_239; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2024 = ret_valid ? _GEN_1490 : dirty_0_240; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2025 = ret_valid ? _GEN_1491 : dirty_0_241; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2026 = ret_valid ? _GEN_1492 : dirty_0_242; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2027 = ret_valid ? _GEN_1493 : dirty_0_243; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2028 = ret_valid ? _GEN_1494 : dirty_0_244; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2029 = ret_valid ? _GEN_1495 : dirty_0_245; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2030 = ret_valid ? _GEN_1496 : dirty_0_246; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2031 = ret_valid ? _GEN_1497 : dirty_0_247; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2032 = ret_valid ? _GEN_1498 : dirty_0_248; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2033 = ret_valid ? _GEN_1499 : dirty_0_249; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2034 = ret_valid ? _GEN_1500 : dirty_0_250; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2035 = ret_valid ? _GEN_1501 : dirty_0_251; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2036 = ret_valid ? _GEN_1502 : dirty_0_252; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2037 = ret_valid ? _GEN_1503 : dirty_0_253; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2038 = ret_valid ? _GEN_1504 : dirty_0_254; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2039 = ret_valid ? _GEN_1505 : dirty_0_255; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2040 = ret_valid ? _GEN_1506 : dirty_1_0; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2041 = ret_valid ? _GEN_1507 : dirty_1_1; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2042 = ret_valid ? _GEN_1508 : dirty_1_2; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2043 = ret_valid ? _GEN_1509 : dirty_1_3; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2044 = ret_valid ? _GEN_1510 : dirty_1_4; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2045 = ret_valid ? _GEN_1511 : dirty_1_5; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2046 = ret_valid ? _GEN_1512 : dirty_1_6; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2047 = ret_valid ? _GEN_1513 : dirty_1_7; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2048 = ret_valid ? _GEN_1514 : dirty_1_8; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2049 = ret_valid ? _GEN_1515 : dirty_1_9; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2050 = ret_valid ? _GEN_1516 : dirty_1_10; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2051 = ret_valid ? _GEN_1517 : dirty_1_11; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2052 = ret_valid ? _GEN_1518 : dirty_1_12; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2053 = ret_valid ? _GEN_1519 : dirty_1_13; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2054 = ret_valid ? _GEN_1520 : dirty_1_14; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2055 = ret_valid ? _GEN_1521 : dirty_1_15; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2056 = ret_valid ? _GEN_1522 : dirty_1_16; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2057 = ret_valid ? _GEN_1523 : dirty_1_17; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2058 = ret_valid ? _GEN_1524 : dirty_1_18; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2059 = ret_valid ? _GEN_1525 : dirty_1_19; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2060 = ret_valid ? _GEN_1526 : dirty_1_20; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2061 = ret_valid ? _GEN_1527 : dirty_1_21; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2062 = ret_valid ? _GEN_1528 : dirty_1_22; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2063 = ret_valid ? _GEN_1529 : dirty_1_23; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2064 = ret_valid ? _GEN_1530 : dirty_1_24; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2065 = ret_valid ? _GEN_1531 : dirty_1_25; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2066 = ret_valid ? _GEN_1532 : dirty_1_26; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2067 = ret_valid ? _GEN_1533 : dirty_1_27; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2068 = ret_valid ? _GEN_1534 : dirty_1_28; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2069 = ret_valid ? _GEN_1535 : dirty_1_29; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2070 = ret_valid ? _GEN_1536 : dirty_1_30; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2071 = ret_valid ? _GEN_1537 : dirty_1_31; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2072 = ret_valid ? _GEN_1538 : dirty_1_32; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2073 = ret_valid ? _GEN_1539 : dirty_1_33; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2074 = ret_valid ? _GEN_1540 : dirty_1_34; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2075 = ret_valid ? _GEN_1541 : dirty_1_35; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2076 = ret_valid ? _GEN_1542 : dirty_1_36; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2077 = ret_valid ? _GEN_1543 : dirty_1_37; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2078 = ret_valid ? _GEN_1544 : dirty_1_38; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2079 = ret_valid ? _GEN_1545 : dirty_1_39; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2080 = ret_valid ? _GEN_1546 : dirty_1_40; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2081 = ret_valid ? _GEN_1547 : dirty_1_41; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2082 = ret_valid ? _GEN_1548 : dirty_1_42; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2083 = ret_valid ? _GEN_1549 : dirty_1_43; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2084 = ret_valid ? _GEN_1550 : dirty_1_44; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2085 = ret_valid ? _GEN_1551 : dirty_1_45; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2086 = ret_valid ? _GEN_1552 : dirty_1_46; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2087 = ret_valid ? _GEN_1553 : dirty_1_47; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2088 = ret_valid ? _GEN_1554 : dirty_1_48; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2089 = ret_valid ? _GEN_1555 : dirty_1_49; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2090 = ret_valid ? _GEN_1556 : dirty_1_50; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2091 = ret_valid ? _GEN_1557 : dirty_1_51; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2092 = ret_valid ? _GEN_1558 : dirty_1_52; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2093 = ret_valid ? _GEN_1559 : dirty_1_53; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2094 = ret_valid ? _GEN_1560 : dirty_1_54; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2095 = ret_valid ? _GEN_1561 : dirty_1_55; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2096 = ret_valid ? _GEN_1562 : dirty_1_56; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2097 = ret_valid ? _GEN_1563 : dirty_1_57; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2098 = ret_valid ? _GEN_1564 : dirty_1_58; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2099 = ret_valid ? _GEN_1565 : dirty_1_59; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2100 = ret_valid ? _GEN_1566 : dirty_1_60; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2101 = ret_valid ? _GEN_1567 : dirty_1_61; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2102 = ret_valid ? _GEN_1568 : dirty_1_62; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2103 = ret_valid ? _GEN_1569 : dirty_1_63; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2104 = ret_valid ? _GEN_1570 : dirty_1_64; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2105 = ret_valid ? _GEN_1571 : dirty_1_65; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2106 = ret_valid ? _GEN_1572 : dirty_1_66; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2107 = ret_valid ? _GEN_1573 : dirty_1_67; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2108 = ret_valid ? _GEN_1574 : dirty_1_68; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2109 = ret_valid ? _GEN_1575 : dirty_1_69; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2110 = ret_valid ? _GEN_1576 : dirty_1_70; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2111 = ret_valid ? _GEN_1577 : dirty_1_71; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2112 = ret_valid ? _GEN_1578 : dirty_1_72; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2113 = ret_valid ? _GEN_1579 : dirty_1_73; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2114 = ret_valid ? _GEN_1580 : dirty_1_74; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2115 = ret_valid ? _GEN_1581 : dirty_1_75; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2116 = ret_valid ? _GEN_1582 : dirty_1_76; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2117 = ret_valid ? _GEN_1583 : dirty_1_77; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2118 = ret_valid ? _GEN_1584 : dirty_1_78; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2119 = ret_valid ? _GEN_1585 : dirty_1_79; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2120 = ret_valid ? _GEN_1586 : dirty_1_80; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2121 = ret_valid ? _GEN_1587 : dirty_1_81; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2122 = ret_valid ? _GEN_1588 : dirty_1_82; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2123 = ret_valid ? _GEN_1589 : dirty_1_83; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2124 = ret_valid ? _GEN_1590 : dirty_1_84; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2125 = ret_valid ? _GEN_1591 : dirty_1_85; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2126 = ret_valid ? _GEN_1592 : dirty_1_86; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2127 = ret_valid ? _GEN_1593 : dirty_1_87; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2128 = ret_valid ? _GEN_1594 : dirty_1_88; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2129 = ret_valid ? _GEN_1595 : dirty_1_89; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2130 = ret_valid ? _GEN_1596 : dirty_1_90; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2131 = ret_valid ? _GEN_1597 : dirty_1_91; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2132 = ret_valid ? _GEN_1598 : dirty_1_92; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2133 = ret_valid ? _GEN_1599 : dirty_1_93; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2134 = ret_valid ? _GEN_1600 : dirty_1_94; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2135 = ret_valid ? _GEN_1601 : dirty_1_95; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2136 = ret_valid ? _GEN_1602 : dirty_1_96; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2137 = ret_valid ? _GEN_1603 : dirty_1_97; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2138 = ret_valid ? _GEN_1604 : dirty_1_98; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2139 = ret_valid ? _GEN_1605 : dirty_1_99; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2140 = ret_valid ? _GEN_1606 : dirty_1_100; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2141 = ret_valid ? _GEN_1607 : dirty_1_101; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2142 = ret_valid ? _GEN_1608 : dirty_1_102; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2143 = ret_valid ? _GEN_1609 : dirty_1_103; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2144 = ret_valid ? _GEN_1610 : dirty_1_104; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2145 = ret_valid ? _GEN_1611 : dirty_1_105; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2146 = ret_valid ? _GEN_1612 : dirty_1_106; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2147 = ret_valid ? _GEN_1613 : dirty_1_107; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2148 = ret_valid ? _GEN_1614 : dirty_1_108; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2149 = ret_valid ? _GEN_1615 : dirty_1_109; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2150 = ret_valid ? _GEN_1616 : dirty_1_110; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2151 = ret_valid ? _GEN_1617 : dirty_1_111; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2152 = ret_valid ? _GEN_1618 : dirty_1_112; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2153 = ret_valid ? _GEN_1619 : dirty_1_113; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2154 = ret_valid ? _GEN_1620 : dirty_1_114; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2155 = ret_valid ? _GEN_1621 : dirty_1_115; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2156 = ret_valid ? _GEN_1622 : dirty_1_116; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2157 = ret_valid ? _GEN_1623 : dirty_1_117; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2158 = ret_valid ? _GEN_1624 : dirty_1_118; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2159 = ret_valid ? _GEN_1625 : dirty_1_119; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2160 = ret_valid ? _GEN_1626 : dirty_1_120; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2161 = ret_valid ? _GEN_1627 : dirty_1_121; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2162 = ret_valid ? _GEN_1628 : dirty_1_122; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2163 = ret_valid ? _GEN_1629 : dirty_1_123; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2164 = ret_valid ? _GEN_1630 : dirty_1_124; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2165 = ret_valid ? _GEN_1631 : dirty_1_125; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2166 = ret_valid ? _GEN_1632 : dirty_1_126; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2167 = ret_valid ? _GEN_1633 : dirty_1_127; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2168 = ret_valid ? _GEN_1634 : dirty_1_128; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2169 = ret_valid ? _GEN_1635 : dirty_1_129; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2170 = ret_valid ? _GEN_1636 : dirty_1_130; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2171 = ret_valid ? _GEN_1637 : dirty_1_131; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2172 = ret_valid ? _GEN_1638 : dirty_1_132; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2173 = ret_valid ? _GEN_1639 : dirty_1_133; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2174 = ret_valid ? _GEN_1640 : dirty_1_134; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2175 = ret_valid ? _GEN_1641 : dirty_1_135; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2176 = ret_valid ? _GEN_1642 : dirty_1_136; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2177 = ret_valid ? _GEN_1643 : dirty_1_137; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2178 = ret_valid ? _GEN_1644 : dirty_1_138; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2179 = ret_valid ? _GEN_1645 : dirty_1_139; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2180 = ret_valid ? _GEN_1646 : dirty_1_140; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2181 = ret_valid ? _GEN_1647 : dirty_1_141; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2182 = ret_valid ? _GEN_1648 : dirty_1_142; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2183 = ret_valid ? _GEN_1649 : dirty_1_143; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2184 = ret_valid ? _GEN_1650 : dirty_1_144; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2185 = ret_valid ? _GEN_1651 : dirty_1_145; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2186 = ret_valid ? _GEN_1652 : dirty_1_146; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2187 = ret_valid ? _GEN_1653 : dirty_1_147; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2188 = ret_valid ? _GEN_1654 : dirty_1_148; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2189 = ret_valid ? _GEN_1655 : dirty_1_149; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2190 = ret_valid ? _GEN_1656 : dirty_1_150; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2191 = ret_valid ? _GEN_1657 : dirty_1_151; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2192 = ret_valid ? _GEN_1658 : dirty_1_152; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2193 = ret_valid ? _GEN_1659 : dirty_1_153; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2194 = ret_valid ? _GEN_1660 : dirty_1_154; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2195 = ret_valid ? _GEN_1661 : dirty_1_155; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2196 = ret_valid ? _GEN_1662 : dirty_1_156; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2197 = ret_valid ? _GEN_1663 : dirty_1_157; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2198 = ret_valid ? _GEN_1664 : dirty_1_158; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2199 = ret_valid ? _GEN_1665 : dirty_1_159; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2200 = ret_valid ? _GEN_1666 : dirty_1_160; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2201 = ret_valid ? _GEN_1667 : dirty_1_161; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2202 = ret_valid ? _GEN_1668 : dirty_1_162; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2203 = ret_valid ? _GEN_1669 : dirty_1_163; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2204 = ret_valid ? _GEN_1670 : dirty_1_164; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2205 = ret_valid ? _GEN_1671 : dirty_1_165; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2206 = ret_valid ? _GEN_1672 : dirty_1_166; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2207 = ret_valid ? _GEN_1673 : dirty_1_167; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2208 = ret_valid ? _GEN_1674 : dirty_1_168; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2209 = ret_valid ? _GEN_1675 : dirty_1_169; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2210 = ret_valid ? _GEN_1676 : dirty_1_170; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2211 = ret_valid ? _GEN_1677 : dirty_1_171; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2212 = ret_valid ? _GEN_1678 : dirty_1_172; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2213 = ret_valid ? _GEN_1679 : dirty_1_173; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2214 = ret_valid ? _GEN_1680 : dirty_1_174; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2215 = ret_valid ? _GEN_1681 : dirty_1_175; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2216 = ret_valid ? _GEN_1682 : dirty_1_176; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2217 = ret_valid ? _GEN_1683 : dirty_1_177; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2218 = ret_valid ? _GEN_1684 : dirty_1_178; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2219 = ret_valid ? _GEN_1685 : dirty_1_179; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2220 = ret_valid ? _GEN_1686 : dirty_1_180; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2221 = ret_valid ? _GEN_1687 : dirty_1_181; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2222 = ret_valid ? _GEN_1688 : dirty_1_182; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2223 = ret_valid ? _GEN_1689 : dirty_1_183; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2224 = ret_valid ? _GEN_1690 : dirty_1_184; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2225 = ret_valid ? _GEN_1691 : dirty_1_185; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2226 = ret_valid ? _GEN_1692 : dirty_1_186; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2227 = ret_valid ? _GEN_1693 : dirty_1_187; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2228 = ret_valid ? _GEN_1694 : dirty_1_188; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2229 = ret_valid ? _GEN_1695 : dirty_1_189; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2230 = ret_valid ? _GEN_1696 : dirty_1_190; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2231 = ret_valid ? _GEN_1697 : dirty_1_191; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2232 = ret_valid ? _GEN_1698 : dirty_1_192; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2233 = ret_valid ? _GEN_1699 : dirty_1_193; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2234 = ret_valid ? _GEN_1700 : dirty_1_194; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2235 = ret_valid ? _GEN_1701 : dirty_1_195; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2236 = ret_valid ? _GEN_1702 : dirty_1_196; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2237 = ret_valid ? _GEN_1703 : dirty_1_197; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2238 = ret_valid ? _GEN_1704 : dirty_1_198; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2239 = ret_valid ? _GEN_1705 : dirty_1_199; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2240 = ret_valid ? _GEN_1706 : dirty_1_200; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2241 = ret_valid ? _GEN_1707 : dirty_1_201; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2242 = ret_valid ? _GEN_1708 : dirty_1_202; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2243 = ret_valid ? _GEN_1709 : dirty_1_203; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2244 = ret_valid ? _GEN_1710 : dirty_1_204; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2245 = ret_valid ? _GEN_1711 : dirty_1_205; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2246 = ret_valid ? _GEN_1712 : dirty_1_206; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2247 = ret_valid ? _GEN_1713 : dirty_1_207; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2248 = ret_valid ? _GEN_1714 : dirty_1_208; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2249 = ret_valid ? _GEN_1715 : dirty_1_209; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2250 = ret_valid ? _GEN_1716 : dirty_1_210; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2251 = ret_valid ? _GEN_1717 : dirty_1_211; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2252 = ret_valid ? _GEN_1718 : dirty_1_212; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2253 = ret_valid ? _GEN_1719 : dirty_1_213; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2254 = ret_valid ? _GEN_1720 : dirty_1_214; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2255 = ret_valid ? _GEN_1721 : dirty_1_215; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2256 = ret_valid ? _GEN_1722 : dirty_1_216; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2257 = ret_valid ? _GEN_1723 : dirty_1_217; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2258 = ret_valid ? _GEN_1724 : dirty_1_218; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2259 = ret_valid ? _GEN_1725 : dirty_1_219; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2260 = ret_valid ? _GEN_1726 : dirty_1_220; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2261 = ret_valid ? _GEN_1727 : dirty_1_221; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2262 = ret_valid ? _GEN_1728 : dirty_1_222; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2263 = ret_valid ? _GEN_1729 : dirty_1_223; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2264 = ret_valid ? _GEN_1730 : dirty_1_224; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2265 = ret_valid ? _GEN_1731 : dirty_1_225; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2266 = ret_valid ? _GEN_1732 : dirty_1_226; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2267 = ret_valid ? _GEN_1733 : dirty_1_227; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2268 = ret_valid ? _GEN_1734 : dirty_1_228; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2269 = ret_valid ? _GEN_1735 : dirty_1_229; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2270 = ret_valid ? _GEN_1736 : dirty_1_230; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2271 = ret_valid ? _GEN_1737 : dirty_1_231; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2272 = ret_valid ? _GEN_1738 : dirty_1_232; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2273 = ret_valid ? _GEN_1739 : dirty_1_233; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2274 = ret_valid ? _GEN_1740 : dirty_1_234; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2275 = ret_valid ? _GEN_1741 : dirty_1_235; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2276 = ret_valid ? _GEN_1742 : dirty_1_236; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2277 = ret_valid ? _GEN_1743 : dirty_1_237; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2278 = ret_valid ? _GEN_1744 : dirty_1_238; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2279 = ret_valid ? _GEN_1745 : dirty_1_239; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2280 = ret_valid ? _GEN_1746 : dirty_1_240; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2281 = ret_valid ? _GEN_1747 : dirty_1_241; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2282 = ret_valid ? _GEN_1748 : dirty_1_242; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2283 = ret_valid ? _GEN_1749 : dirty_1_243; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2284 = ret_valid ? _GEN_1750 : dirty_1_244; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2285 = ret_valid ? _GEN_1751 : dirty_1_245; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2286 = ret_valid ? _GEN_1752 : dirty_1_246; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2287 = ret_valid ? _GEN_1753 : dirty_1_247; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2288 = ret_valid ? _GEN_1754 : dirty_1_248; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2289 = ret_valid ? _GEN_1755 : dirty_1_249; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2290 = ret_valid ? _GEN_1756 : dirty_1_250; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2291 = ret_valid ? _GEN_1757 : dirty_1_251; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2292 = ret_valid ? _GEN_1758 : dirty_1_252; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2293 = ret_valid ? _GEN_1759 : dirty_1_253; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2294 = ret_valid ? _GEN_1760 : dirty_1_254; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2295 = ret_valid ? _GEN_1761 : dirty_1_255; // @[dcache.scala 384:17 113:28]
  wire  _GEN_2296 = ret_valid & _GEN_1762; // @[dcache.scala 384:17 144:25]
  wire  _GEN_2297 = ret_valid & _GEN_1763; // @[dcache.scala 384:17 144:25]
  wire [20:0] _GEN_2298 = ret_valid ? _GEN_1764 : 21'h0; // @[dcache.scala 384:17 143:25]
  wire [20:0] _GEN_2299 = ret_valid ? _GEN_1765 : 21'h0; // @[dcache.scala 384:17 143:25]
  wire  _T_51 = ret_valid & ret_last; // @[dcache.scala 398:32]
  wire [31:0] _GEN_2301 = _T_51 ? ret_data : 32'h7777; // @[dcache.scala 399:17 155:25 401:61]
  wire [2:0] _GEN_2302 = _T_51 ? 3'h0 : 3'h5; // @[dcache.scala 399:17 380:41 402:61]
  wire  _GEN_2303 = _T_51 ? 1'h0 : req_valid; // @[dcache.scala 399:17 116:34 403:61]
  wire [20:0] _GEN_2305 = waySel ? tagv_r_1 : tagv_r_0; // @[dcache.scala 409:{106,106}]
  wire  _GEN_13518 = ~waySel; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2307 = ~waySel & _GEN_11959 ? dirty_0_1 : dirty_0_0; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2308 = ~waySel & _GEN_11961 ? dirty_0_2 : _GEN_2307; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2309 = ~waySel & _GEN_11963 ? dirty_0_3 : _GEN_2308; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2310 = ~waySel & _GEN_11965 ? dirty_0_4 : _GEN_2309; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2311 = ~waySel & _GEN_11967 ? dirty_0_5 : _GEN_2310; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2312 = ~waySel & _GEN_11969 ? dirty_0_6 : _GEN_2311; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2313 = ~waySel & _GEN_11971 ? dirty_0_7 : _GEN_2312; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2314 = ~waySel & _GEN_11973 ? dirty_0_8 : _GEN_2313; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2315 = ~waySel & _GEN_11975 ? dirty_0_9 : _GEN_2314; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2316 = ~waySel & _GEN_11977 ? dirty_0_10 : _GEN_2315; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2317 = ~waySel & _GEN_11979 ? dirty_0_11 : _GEN_2316; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2318 = ~waySel & _GEN_11981 ? dirty_0_12 : _GEN_2317; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2319 = ~waySel & _GEN_11983 ? dirty_0_13 : _GEN_2318; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2320 = ~waySel & _GEN_11985 ? dirty_0_14 : _GEN_2319; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2321 = ~waySel & _GEN_11987 ? dirty_0_15 : _GEN_2320; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2322 = ~waySel & _GEN_11989 ? dirty_0_16 : _GEN_2321; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2323 = ~waySel & _GEN_11991 ? dirty_0_17 : _GEN_2322; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2324 = ~waySel & _GEN_11993 ? dirty_0_18 : _GEN_2323; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2325 = ~waySel & _GEN_11995 ? dirty_0_19 : _GEN_2324; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2326 = ~waySel & _GEN_11997 ? dirty_0_20 : _GEN_2325; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2327 = ~waySel & _GEN_11999 ? dirty_0_21 : _GEN_2326; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2328 = ~waySel & _GEN_12001 ? dirty_0_22 : _GEN_2327; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2329 = ~waySel & _GEN_12003 ? dirty_0_23 : _GEN_2328; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2330 = ~waySel & _GEN_12005 ? dirty_0_24 : _GEN_2329; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2331 = ~waySel & _GEN_12007 ? dirty_0_25 : _GEN_2330; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2332 = ~waySel & _GEN_12009 ? dirty_0_26 : _GEN_2331; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2333 = ~waySel & _GEN_12011 ? dirty_0_27 : _GEN_2332; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2334 = ~waySel & _GEN_12013 ? dirty_0_28 : _GEN_2333; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2335 = ~waySel & _GEN_12015 ? dirty_0_29 : _GEN_2334; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2336 = ~waySel & _GEN_12017 ? dirty_0_30 : _GEN_2335; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2337 = ~waySel & _GEN_12019 ? dirty_0_31 : _GEN_2336; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2338 = ~waySel & _GEN_12021 ? dirty_0_32 : _GEN_2337; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2339 = ~waySel & _GEN_12023 ? dirty_0_33 : _GEN_2338; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2340 = ~waySel & _GEN_12025 ? dirty_0_34 : _GEN_2339; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2341 = ~waySel & _GEN_12027 ? dirty_0_35 : _GEN_2340; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2342 = ~waySel & _GEN_12029 ? dirty_0_36 : _GEN_2341; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2343 = ~waySel & _GEN_12031 ? dirty_0_37 : _GEN_2342; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2344 = ~waySel & _GEN_12033 ? dirty_0_38 : _GEN_2343; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2345 = ~waySel & _GEN_12035 ? dirty_0_39 : _GEN_2344; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2346 = ~waySel & _GEN_12037 ? dirty_0_40 : _GEN_2345; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2347 = ~waySel & _GEN_12039 ? dirty_0_41 : _GEN_2346; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2348 = ~waySel & _GEN_12041 ? dirty_0_42 : _GEN_2347; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2349 = ~waySel & _GEN_12043 ? dirty_0_43 : _GEN_2348; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2350 = ~waySel & _GEN_12045 ? dirty_0_44 : _GEN_2349; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2351 = ~waySel & _GEN_12047 ? dirty_0_45 : _GEN_2350; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2352 = ~waySel & _GEN_12049 ? dirty_0_46 : _GEN_2351; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2353 = ~waySel & _GEN_12051 ? dirty_0_47 : _GEN_2352; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2354 = ~waySel & _GEN_12053 ? dirty_0_48 : _GEN_2353; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2355 = ~waySel & _GEN_12055 ? dirty_0_49 : _GEN_2354; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2356 = ~waySel & _GEN_12057 ? dirty_0_50 : _GEN_2355; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2357 = ~waySel & _GEN_12059 ? dirty_0_51 : _GEN_2356; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2358 = ~waySel & _GEN_12061 ? dirty_0_52 : _GEN_2357; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2359 = ~waySel & _GEN_12063 ? dirty_0_53 : _GEN_2358; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2360 = ~waySel & _GEN_12065 ? dirty_0_54 : _GEN_2359; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2361 = ~waySel & _GEN_12067 ? dirty_0_55 : _GEN_2360; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2362 = ~waySel & _GEN_12069 ? dirty_0_56 : _GEN_2361; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2363 = ~waySel & _GEN_12071 ? dirty_0_57 : _GEN_2362; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2364 = ~waySel & _GEN_12073 ? dirty_0_58 : _GEN_2363; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2365 = ~waySel & _GEN_12075 ? dirty_0_59 : _GEN_2364; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2366 = ~waySel & _GEN_12077 ? dirty_0_60 : _GEN_2365; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2367 = ~waySel & _GEN_12079 ? dirty_0_61 : _GEN_2366; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2368 = ~waySel & _GEN_12081 ? dirty_0_62 : _GEN_2367; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2369 = ~waySel & _GEN_12083 ? dirty_0_63 : _GEN_2368; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2370 = ~waySel & _GEN_12085 ? dirty_0_64 : _GEN_2369; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2371 = ~waySel & _GEN_12087 ? dirty_0_65 : _GEN_2370; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2372 = ~waySel & _GEN_12089 ? dirty_0_66 : _GEN_2371; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2373 = ~waySel & _GEN_12091 ? dirty_0_67 : _GEN_2372; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2374 = ~waySel & _GEN_12093 ? dirty_0_68 : _GEN_2373; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2375 = ~waySel & _GEN_12095 ? dirty_0_69 : _GEN_2374; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2376 = ~waySel & _GEN_12097 ? dirty_0_70 : _GEN_2375; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2377 = ~waySel & _GEN_12099 ? dirty_0_71 : _GEN_2376; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2378 = ~waySel & _GEN_12101 ? dirty_0_72 : _GEN_2377; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2379 = ~waySel & _GEN_12103 ? dirty_0_73 : _GEN_2378; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2380 = ~waySel & _GEN_12105 ? dirty_0_74 : _GEN_2379; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2381 = ~waySel & _GEN_12107 ? dirty_0_75 : _GEN_2380; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2382 = ~waySel & _GEN_12109 ? dirty_0_76 : _GEN_2381; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2383 = ~waySel & _GEN_12111 ? dirty_0_77 : _GEN_2382; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2384 = ~waySel & _GEN_12113 ? dirty_0_78 : _GEN_2383; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2385 = ~waySel & _GEN_12115 ? dirty_0_79 : _GEN_2384; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2386 = ~waySel & _GEN_12117 ? dirty_0_80 : _GEN_2385; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2387 = ~waySel & _GEN_12119 ? dirty_0_81 : _GEN_2386; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2388 = ~waySel & _GEN_12121 ? dirty_0_82 : _GEN_2387; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2389 = ~waySel & _GEN_12123 ? dirty_0_83 : _GEN_2388; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2390 = ~waySel & _GEN_12125 ? dirty_0_84 : _GEN_2389; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2391 = ~waySel & _GEN_12127 ? dirty_0_85 : _GEN_2390; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2392 = ~waySel & _GEN_12129 ? dirty_0_86 : _GEN_2391; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2393 = ~waySel & _GEN_12131 ? dirty_0_87 : _GEN_2392; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2394 = ~waySel & _GEN_12133 ? dirty_0_88 : _GEN_2393; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2395 = ~waySel & _GEN_12135 ? dirty_0_89 : _GEN_2394; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2396 = ~waySel & _GEN_12137 ? dirty_0_90 : _GEN_2395; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2397 = ~waySel & _GEN_12139 ? dirty_0_91 : _GEN_2396; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2398 = ~waySel & _GEN_12141 ? dirty_0_92 : _GEN_2397; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2399 = ~waySel & _GEN_12143 ? dirty_0_93 : _GEN_2398; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2400 = ~waySel & _GEN_12145 ? dirty_0_94 : _GEN_2399; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2401 = ~waySel & _GEN_12147 ? dirty_0_95 : _GEN_2400; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2402 = ~waySel & _GEN_12149 ? dirty_0_96 : _GEN_2401; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2403 = ~waySel & _GEN_12151 ? dirty_0_97 : _GEN_2402; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2404 = ~waySel & _GEN_12153 ? dirty_0_98 : _GEN_2403; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2405 = ~waySel & _GEN_12155 ? dirty_0_99 : _GEN_2404; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2406 = ~waySel & _GEN_12157 ? dirty_0_100 : _GEN_2405; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2407 = ~waySel & _GEN_12159 ? dirty_0_101 : _GEN_2406; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2408 = ~waySel & _GEN_12161 ? dirty_0_102 : _GEN_2407; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2409 = ~waySel & _GEN_12163 ? dirty_0_103 : _GEN_2408; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2410 = ~waySel & _GEN_12165 ? dirty_0_104 : _GEN_2409; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2411 = ~waySel & _GEN_12167 ? dirty_0_105 : _GEN_2410; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2412 = ~waySel & _GEN_12169 ? dirty_0_106 : _GEN_2411; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2413 = ~waySel & _GEN_12171 ? dirty_0_107 : _GEN_2412; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2414 = ~waySel & _GEN_12173 ? dirty_0_108 : _GEN_2413; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2415 = ~waySel & _GEN_12175 ? dirty_0_109 : _GEN_2414; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2416 = ~waySel & _GEN_12177 ? dirty_0_110 : _GEN_2415; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2417 = ~waySel & _GEN_12179 ? dirty_0_111 : _GEN_2416; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2418 = ~waySel & _GEN_12181 ? dirty_0_112 : _GEN_2417; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2419 = ~waySel & _GEN_12183 ? dirty_0_113 : _GEN_2418; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2420 = ~waySel & _GEN_12185 ? dirty_0_114 : _GEN_2419; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2421 = ~waySel & _GEN_12187 ? dirty_0_115 : _GEN_2420; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2422 = ~waySel & _GEN_12189 ? dirty_0_116 : _GEN_2421; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2423 = ~waySel & _GEN_12191 ? dirty_0_117 : _GEN_2422; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2424 = ~waySel & _GEN_12193 ? dirty_0_118 : _GEN_2423; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2425 = ~waySel & _GEN_12195 ? dirty_0_119 : _GEN_2424; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2426 = ~waySel & _GEN_12197 ? dirty_0_120 : _GEN_2425; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2427 = ~waySel & _GEN_12199 ? dirty_0_121 : _GEN_2426; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2428 = ~waySel & _GEN_12201 ? dirty_0_122 : _GEN_2427; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2429 = ~waySel & _GEN_12203 ? dirty_0_123 : _GEN_2428; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2430 = ~waySel & _GEN_12205 ? dirty_0_124 : _GEN_2429; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2431 = ~waySel & _GEN_12207 ? dirty_0_125 : _GEN_2430; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2432 = ~waySel & _GEN_12209 ? dirty_0_126 : _GEN_2431; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2433 = ~waySel & _GEN_12211 ? dirty_0_127 : _GEN_2432; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2434 = ~waySel & _GEN_12213 ? dirty_0_128 : _GEN_2433; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2435 = ~waySel & _GEN_12215 ? dirty_0_129 : _GEN_2434; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2436 = ~waySel & _GEN_12217 ? dirty_0_130 : _GEN_2435; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2437 = ~waySel & _GEN_12219 ? dirty_0_131 : _GEN_2436; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2438 = ~waySel & _GEN_12221 ? dirty_0_132 : _GEN_2437; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2439 = ~waySel & _GEN_12223 ? dirty_0_133 : _GEN_2438; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2440 = ~waySel & _GEN_12225 ? dirty_0_134 : _GEN_2439; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2441 = ~waySel & _GEN_12227 ? dirty_0_135 : _GEN_2440; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2442 = ~waySel & _GEN_12229 ? dirty_0_136 : _GEN_2441; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2443 = ~waySel & _GEN_12231 ? dirty_0_137 : _GEN_2442; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2444 = ~waySel & _GEN_12233 ? dirty_0_138 : _GEN_2443; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2445 = ~waySel & _GEN_12235 ? dirty_0_139 : _GEN_2444; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2446 = ~waySel & _GEN_12237 ? dirty_0_140 : _GEN_2445; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2447 = ~waySel & _GEN_12239 ? dirty_0_141 : _GEN_2446; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2448 = ~waySel & _GEN_12241 ? dirty_0_142 : _GEN_2447; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2449 = ~waySel & _GEN_12243 ? dirty_0_143 : _GEN_2448; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2450 = ~waySel & _GEN_12245 ? dirty_0_144 : _GEN_2449; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2451 = ~waySel & _GEN_12247 ? dirty_0_145 : _GEN_2450; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2452 = ~waySel & _GEN_12249 ? dirty_0_146 : _GEN_2451; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2453 = ~waySel & _GEN_12251 ? dirty_0_147 : _GEN_2452; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2454 = ~waySel & _GEN_12253 ? dirty_0_148 : _GEN_2453; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2455 = ~waySel & _GEN_12255 ? dirty_0_149 : _GEN_2454; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2456 = ~waySel & _GEN_12257 ? dirty_0_150 : _GEN_2455; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2457 = ~waySel & _GEN_12259 ? dirty_0_151 : _GEN_2456; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2458 = ~waySel & _GEN_12261 ? dirty_0_152 : _GEN_2457; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2459 = ~waySel & _GEN_12263 ? dirty_0_153 : _GEN_2458; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2460 = ~waySel & _GEN_12265 ? dirty_0_154 : _GEN_2459; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2461 = ~waySel & _GEN_12267 ? dirty_0_155 : _GEN_2460; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2462 = ~waySel & _GEN_12269 ? dirty_0_156 : _GEN_2461; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2463 = ~waySel & _GEN_12271 ? dirty_0_157 : _GEN_2462; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2464 = ~waySel & _GEN_12273 ? dirty_0_158 : _GEN_2463; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2465 = ~waySel & _GEN_12275 ? dirty_0_159 : _GEN_2464; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2466 = ~waySel & _GEN_12277 ? dirty_0_160 : _GEN_2465; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2467 = ~waySel & _GEN_12279 ? dirty_0_161 : _GEN_2466; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2468 = ~waySel & _GEN_12281 ? dirty_0_162 : _GEN_2467; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2469 = ~waySel & _GEN_12283 ? dirty_0_163 : _GEN_2468; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2470 = ~waySel & _GEN_12285 ? dirty_0_164 : _GEN_2469; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2471 = ~waySel & _GEN_12287 ? dirty_0_165 : _GEN_2470; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2472 = ~waySel & _GEN_12289 ? dirty_0_166 : _GEN_2471; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2473 = ~waySel & _GEN_12291 ? dirty_0_167 : _GEN_2472; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2474 = ~waySel & _GEN_12293 ? dirty_0_168 : _GEN_2473; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2475 = ~waySel & _GEN_12295 ? dirty_0_169 : _GEN_2474; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2476 = ~waySel & _GEN_12297 ? dirty_0_170 : _GEN_2475; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2477 = ~waySel & _GEN_12299 ? dirty_0_171 : _GEN_2476; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2478 = ~waySel & _GEN_12301 ? dirty_0_172 : _GEN_2477; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2479 = ~waySel & _GEN_12303 ? dirty_0_173 : _GEN_2478; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2480 = ~waySel & _GEN_12305 ? dirty_0_174 : _GEN_2479; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2481 = ~waySel & _GEN_12307 ? dirty_0_175 : _GEN_2480; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2482 = ~waySel & _GEN_12309 ? dirty_0_176 : _GEN_2481; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2483 = ~waySel & _GEN_12311 ? dirty_0_177 : _GEN_2482; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2484 = ~waySel & _GEN_12313 ? dirty_0_178 : _GEN_2483; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2485 = ~waySel & _GEN_12315 ? dirty_0_179 : _GEN_2484; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2486 = ~waySel & _GEN_12317 ? dirty_0_180 : _GEN_2485; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2487 = ~waySel & _GEN_12319 ? dirty_0_181 : _GEN_2486; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2488 = ~waySel & _GEN_12321 ? dirty_0_182 : _GEN_2487; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2489 = ~waySel & _GEN_12323 ? dirty_0_183 : _GEN_2488; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2490 = ~waySel & _GEN_12325 ? dirty_0_184 : _GEN_2489; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2491 = ~waySel & _GEN_12327 ? dirty_0_185 : _GEN_2490; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2492 = ~waySel & _GEN_12329 ? dirty_0_186 : _GEN_2491; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2493 = ~waySel & _GEN_12331 ? dirty_0_187 : _GEN_2492; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2494 = ~waySel & _GEN_12333 ? dirty_0_188 : _GEN_2493; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2495 = ~waySel & _GEN_12335 ? dirty_0_189 : _GEN_2494; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2496 = ~waySel & _GEN_12337 ? dirty_0_190 : _GEN_2495; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2497 = ~waySel & _GEN_12339 ? dirty_0_191 : _GEN_2496; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2498 = ~waySel & _GEN_12341 ? dirty_0_192 : _GEN_2497; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2499 = ~waySel & _GEN_12343 ? dirty_0_193 : _GEN_2498; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2500 = ~waySel & _GEN_12345 ? dirty_0_194 : _GEN_2499; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2501 = ~waySel & _GEN_12347 ? dirty_0_195 : _GEN_2500; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2502 = ~waySel & _GEN_12349 ? dirty_0_196 : _GEN_2501; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2503 = ~waySel & _GEN_12351 ? dirty_0_197 : _GEN_2502; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2504 = ~waySel & _GEN_12353 ? dirty_0_198 : _GEN_2503; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2505 = ~waySel & _GEN_12355 ? dirty_0_199 : _GEN_2504; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2506 = ~waySel & _GEN_12357 ? dirty_0_200 : _GEN_2505; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2507 = ~waySel & _GEN_12359 ? dirty_0_201 : _GEN_2506; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2508 = ~waySel & _GEN_12361 ? dirty_0_202 : _GEN_2507; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2509 = ~waySel & _GEN_12363 ? dirty_0_203 : _GEN_2508; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2510 = ~waySel & _GEN_12365 ? dirty_0_204 : _GEN_2509; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2511 = ~waySel & _GEN_12367 ? dirty_0_205 : _GEN_2510; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2512 = ~waySel & _GEN_12369 ? dirty_0_206 : _GEN_2511; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2513 = ~waySel & _GEN_12371 ? dirty_0_207 : _GEN_2512; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2514 = ~waySel & _GEN_12373 ? dirty_0_208 : _GEN_2513; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2515 = ~waySel & _GEN_12375 ? dirty_0_209 : _GEN_2514; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2516 = ~waySel & _GEN_12377 ? dirty_0_210 : _GEN_2515; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2517 = ~waySel & _GEN_12379 ? dirty_0_211 : _GEN_2516; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2518 = ~waySel & _GEN_12381 ? dirty_0_212 : _GEN_2517; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2519 = ~waySel & _GEN_12383 ? dirty_0_213 : _GEN_2518; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2520 = ~waySel & _GEN_12385 ? dirty_0_214 : _GEN_2519; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2521 = ~waySel & _GEN_12387 ? dirty_0_215 : _GEN_2520; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2522 = ~waySel & _GEN_12389 ? dirty_0_216 : _GEN_2521; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2523 = ~waySel & _GEN_12391 ? dirty_0_217 : _GEN_2522; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2524 = ~waySel & _GEN_12393 ? dirty_0_218 : _GEN_2523; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2525 = ~waySel & _GEN_12395 ? dirty_0_219 : _GEN_2524; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2526 = ~waySel & _GEN_12397 ? dirty_0_220 : _GEN_2525; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2527 = ~waySel & _GEN_12399 ? dirty_0_221 : _GEN_2526; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2528 = ~waySel & _GEN_12401 ? dirty_0_222 : _GEN_2527; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2529 = ~waySel & _GEN_12403 ? dirty_0_223 : _GEN_2528; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2530 = ~waySel & _GEN_12405 ? dirty_0_224 : _GEN_2529; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2531 = ~waySel & _GEN_12407 ? dirty_0_225 : _GEN_2530; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2532 = ~waySel & _GEN_12409 ? dirty_0_226 : _GEN_2531; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2533 = ~waySel & _GEN_12411 ? dirty_0_227 : _GEN_2532; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2534 = ~waySel & _GEN_12413 ? dirty_0_228 : _GEN_2533; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2535 = ~waySel & _GEN_12415 ? dirty_0_229 : _GEN_2534; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2536 = ~waySel & _GEN_12417 ? dirty_0_230 : _GEN_2535; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2537 = ~waySel & _GEN_12419 ? dirty_0_231 : _GEN_2536; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2538 = ~waySel & _GEN_12421 ? dirty_0_232 : _GEN_2537; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2539 = ~waySel & _GEN_12423 ? dirty_0_233 : _GEN_2538; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2540 = ~waySel & _GEN_12425 ? dirty_0_234 : _GEN_2539; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2541 = ~waySel & _GEN_12427 ? dirty_0_235 : _GEN_2540; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2542 = ~waySel & _GEN_12429 ? dirty_0_236 : _GEN_2541; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2543 = ~waySel & _GEN_12431 ? dirty_0_237 : _GEN_2542; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2544 = ~waySel & _GEN_12433 ? dirty_0_238 : _GEN_2543; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2545 = ~waySel & _GEN_12435 ? dirty_0_239 : _GEN_2544; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2546 = ~waySel & _GEN_12437 ? dirty_0_240 : _GEN_2545; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2547 = ~waySel & _GEN_12439 ? dirty_0_241 : _GEN_2546; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2548 = ~waySel & _GEN_12441 ? dirty_0_242 : _GEN_2547; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2549 = ~waySel & _GEN_12443 ? dirty_0_243 : _GEN_2548; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2550 = ~waySel & _GEN_12445 ? dirty_0_244 : _GEN_2549; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2551 = ~waySel & _GEN_12447 ? dirty_0_245 : _GEN_2550; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2552 = ~waySel & _GEN_12449 ? dirty_0_246 : _GEN_2551; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2553 = ~waySel & _GEN_12451 ? dirty_0_247 : _GEN_2552; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2554 = ~waySel & _GEN_12453 ? dirty_0_248 : _GEN_2553; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2555 = ~waySel & _GEN_12455 ? dirty_0_249 : _GEN_2554; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2556 = ~waySel & _GEN_12457 ? dirty_0_250 : _GEN_2555; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2557 = ~waySel & _GEN_12459 ? dirty_0_251 : _GEN_2556; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2558 = ~waySel & _GEN_12461 ? dirty_0_252 : _GEN_2557; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2559 = ~waySel & _GEN_12463 ? dirty_0_253 : _GEN_2558; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2560 = ~waySel & _GEN_12465 ? dirty_0_254 : _GEN_2559; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2561 = ~waySel & _GEN_12467 ? dirty_0_255 : _GEN_2560; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2562 = waySel & _GEN_12468 ? dirty_1_0 : _GEN_2561; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2563 = waySel & _GEN_11959 ? dirty_1_1 : _GEN_2562; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2564 = waySel & _GEN_11961 ? dirty_1_2 : _GEN_2563; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2565 = waySel & _GEN_11963 ? dirty_1_3 : _GEN_2564; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2566 = waySel & _GEN_11965 ? dirty_1_4 : _GEN_2565; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2567 = waySel & _GEN_11967 ? dirty_1_5 : _GEN_2566; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2568 = waySel & _GEN_11969 ? dirty_1_6 : _GEN_2567; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2569 = waySel & _GEN_11971 ? dirty_1_7 : _GEN_2568; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2570 = waySel & _GEN_11973 ? dirty_1_8 : _GEN_2569; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2571 = waySel & _GEN_11975 ? dirty_1_9 : _GEN_2570; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2572 = waySel & _GEN_11977 ? dirty_1_10 : _GEN_2571; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2573 = waySel & _GEN_11979 ? dirty_1_11 : _GEN_2572; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2574 = waySel & _GEN_11981 ? dirty_1_12 : _GEN_2573; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2575 = waySel & _GEN_11983 ? dirty_1_13 : _GEN_2574; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2576 = waySel & _GEN_11985 ? dirty_1_14 : _GEN_2575; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2577 = waySel & _GEN_11987 ? dirty_1_15 : _GEN_2576; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2578 = waySel & _GEN_11989 ? dirty_1_16 : _GEN_2577; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2579 = waySel & _GEN_11991 ? dirty_1_17 : _GEN_2578; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2580 = waySel & _GEN_11993 ? dirty_1_18 : _GEN_2579; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2581 = waySel & _GEN_11995 ? dirty_1_19 : _GEN_2580; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2582 = waySel & _GEN_11997 ? dirty_1_20 : _GEN_2581; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2583 = waySel & _GEN_11999 ? dirty_1_21 : _GEN_2582; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2584 = waySel & _GEN_12001 ? dirty_1_22 : _GEN_2583; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2585 = waySel & _GEN_12003 ? dirty_1_23 : _GEN_2584; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2586 = waySel & _GEN_12005 ? dirty_1_24 : _GEN_2585; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2587 = waySel & _GEN_12007 ? dirty_1_25 : _GEN_2586; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2588 = waySel & _GEN_12009 ? dirty_1_26 : _GEN_2587; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2589 = waySel & _GEN_12011 ? dirty_1_27 : _GEN_2588; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2590 = waySel & _GEN_12013 ? dirty_1_28 : _GEN_2589; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2591 = waySel & _GEN_12015 ? dirty_1_29 : _GEN_2590; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2592 = waySel & _GEN_12017 ? dirty_1_30 : _GEN_2591; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2593 = waySel & _GEN_12019 ? dirty_1_31 : _GEN_2592; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2594 = waySel & _GEN_12021 ? dirty_1_32 : _GEN_2593; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2595 = waySel & _GEN_12023 ? dirty_1_33 : _GEN_2594; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2596 = waySel & _GEN_12025 ? dirty_1_34 : _GEN_2595; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2597 = waySel & _GEN_12027 ? dirty_1_35 : _GEN_2596; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2598 = waySel & _GEN_12029 ? dirty_1_36 : _GEN_2597; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2599 = waySel & _GEN_12031 ? dirty_1_37 : _GEN_2598; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2600 = waySel & _GEN_12033 ? dirty_1_38 : _GEN_2599; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2601 = waySel & _GEN_12035 ? dirty_1_39 : _GEN_2600; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2602 = waySel & _GEN_12037 ? dirty_1_40 : _GEN_2601; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2603 = waySel & _GEN_12039 ? dirty_1_41 : _GEN_2602; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2604 = waySel & _GEN_12041 ? dirty_1_42 : _GEN_2603; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2605 = waySel & _GEN_12043 ? dirty_1_43 : _GEN_2604; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2606 = waySel & _GEN_12045 ? dirty_1_44 : _GEN_2605; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2607 = waySel & _GEN_12047 ? dirty_1_45 : _GEN_2606; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2608 = waySel & _GEN_12049 ? dirty_1_46 : _GEN_2607; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2609 = waySel & _GEN_12051 ? dirty_1_47 : _GEN_2608; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2610 = waySel & _GEN_12053 ? dirty_1_48 : _GEN_2609; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2611 = waySel & _GEN_12055 ? dirty_1_49 : _GEN_2610; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2612 = waySel & _GEN_12057 ? dirty_1_50 : _GEN_2611; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2613 = waySel & _GEN_12059 ? dirty_1_51 : _GEN_2612; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2614 = waySel & _GEN_12061 ? dirty_1_52 : _GEN_2613; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2615 = waySel & _GEN_12063 ? dirty_1_53 : _GEN_2614; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2616 = waySel & _GEN_12065 ? dirty_1_54 : _GEN_2615; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2617 = waySel & _GEN_12067 ? dirty_1_55 : _GEN_2616; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2618 = waySel & _GEN_12069 ? dirty_1_56 : _GEN_2617; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2619 = waySel & _GEN_12071 ? dirty_1_57 : _GEN_2618; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2620 = waySel & _GEN_12073 ? dirty_1_58 : _GEN_2619; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2621 = waySel & _GEN_12075 ? dirty_1_59 : _GEN_2620; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2622 = waySel & _GEN_12077 ? dirty_1_60 : _GEN_2621; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2623 = waySel & _GEN_12079 ? dirty_1_61 : _GEN_2622; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2624 = waySel & _GEN_12081 ? dirty_1_62 : _GEN_2623; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2625 = waySel & _GEN_12083 ? dirty_1_63 : _GEN_2624; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2626 = waySel & _GEN_12085 ? dirty_1_64 : _GEN_2625; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2627 = waySel & _GEN_12087 ? dirty_1_65 : _GEN_2626; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2628 = waySel & _GEN_12089 ? dirty_1_66 : _GEN_2627; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2629 = waySel & _GEN_12091 ? dirty_1_67 : _GEN_2628; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2630 = waySel & _GEN_12093 ? dirty_1_68 : _GEN_2629; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2631 = waySel & _GEN_12095 ? dirty_1_69 : _GEN_2630; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2632 = waySel & _GEN_12097 ? dirty_1_70 : _GEN_2631; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2633 = waySel & _GEN_12099 ? dirty_1_71 : _GEN_2632; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2634 = waySel & _GEN_12101 ? dirty_1_72 : _GEN_2633; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2635 = waySel & _GEN_12103 ? dirty_1_73 : _GEN_2634; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2636 = waySel & _GEN_12105 ? dirty_1_74 : _GEN_2635; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2637 = waySel & _GEN_12107 ? dirty_1_75 : _GEN_2636; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2638 = waySel & _GEN_12109 ? dirty_1_76 : _GEN_2637; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2639 = waySel & _GEN_12111 ? dirty_1_77 : _GEN_2638; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2640 = waySel & _GEN_12113 ? dirty_1_78 : _GEN_2639; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2641 = waySel & _GEN_12115 ? dirty_1_79 : _GEN_2640; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2642 = waySel & _GEN_12117 ? dirty_1_80 : _GEN_2641; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2643 = waySel & _GEN_12119 ? dirty_1_81 : _GEN_2642; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2644 = waySel & _GEN_12121 ? dirty_1_82 : _GEN_2643; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2645 = waySel & _GEN_12123 ? dirty_1_83 : _GEN_2644; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2646 = waySel & _GEN_12125 ? dirty_1_84 : _GEN_2645; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2647 = waySel & _GEN_12127 ? dirty_1_85 : _GEN_2646; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2648 = waySel & _GEN_12129 ? dirty_1_86 : _GEN_2647; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2649 = waySel & _GEN_12131 ? dirty_1_87 : _GEN_2648; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2650 = waySel & _GEN_12133 ? dirty_1_88 : _GEN_2649; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2651 = waySel & _GEN_12135 ? dirty_1_89 : _GEN_2650; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2652 = waySel & _GEN_12137 ? dirty_1_90 : _GEN_2651; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2653 = waySel & _GEN_12139 ? dirty_1_91 : _GEN_2652; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2654 = waySel & _GEN_12141 ? dirty_1_92 : _GEN_2653; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2655 = waySel & _GEN_12143 ? dirty_1_93 : _GEN_2654; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2656 = waySel & _GEN_12145 ? dirty_1_94 : _GEN_2655; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2657 = waySel & _GEN_12147 ? dirty_1_95 : _GEN_2656; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2658 = waySel & _GEN_12149 ? dirty_1_96 : _GEN_2657; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2659 = waySel & _GEN_12151 ? dirty_1_97 : _GEN_2658; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2660 = waySel & _GEN_12153 ? dirty_1_98 : _GEN_2659; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2661 = waySel & _GEN_12155 ? dirty_1_99 : _GEN_2660; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2662 = waySel & _GEN_12157 ? dirty_1_100 : _GEN_2661; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2663 = waySel & _GEN_12159 ? dirty_1_101 : _GEN_2662; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2664 = waySel & _GEN_12161 ? dirty_1_102 : _GEN_2663; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2665 = waySel & _GEN_12163 ? dirty_1_103 : _GEN_2664; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2666 = waySel & _GEN_12165 ? dirty_1_104 : _GEN_2665; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2667 = waySel & _GEN_12167 ? dirty_1_105 : _GEN_2666; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2668 = waySel & _GEN_12169 ? dirty_1_106 : _GEN_2667; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2669 = waySel & _GEN_12171 ? dirty_1_107 : _GEN_2668; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2670 = waySel & _GEN_12173 ? dirty_1_108 : _GEN_2669; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2671 = waySel & _GEN_12175 ? dirty_1_109 : _GEN_2670; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2672 = waySel & _GEN_12177 ? dirty_1_110 : _GEN_2671; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2673 = waySel & _GEN_12179 ? dirty_1_111 : _GEN_2672; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2674 = waySel & _GEN_12181 ? dirty_1_112 : _GEN_2673; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2675 = waySel & _GEN_12183 ? dirty_1_113 : _GEN_2674; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2676 = waySel & _GEN_12185 ? dirty_1_114 : _GEN_2675; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2677 = waySel & _GEN_12187 ? dirty_1_115 : _GEN_2676; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2678 = waySel & _GEN_12189 ? dirty_1_116 : _GEN_2677; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2679 = waySel & _GEN_12191 ? dirty_1_117 : _GEN_2678; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2680 = waySel & _GEN_12193 ? dirty_1_118 : _GEN_2679; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2681 = waySel & _GEN_12195 ? dirty_1_119 : _GEN_2680; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2682 = waySel & _GEN_12197 ? dirty_1_120 : _GEN_2681; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2683 = waySel & _GEN_12199 ? dirty_1_121 : _GEN_2682; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2684 = waySel & _GEN_12201 ? dirty_1_122 : _GEN_2683; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2685 = waySel & _GEN_12203 ? dirty_1_123 : _GEN_2684; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2686 = waySel & _GEN_12205 ? dirty_1_124 : _GEN_2685; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2687 = waySel & _GEN_12207 ? dirty_1_125 : _GEN_2686; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2688 = waySel & _GEN_12209 ? dirty_1_126 : _GEN_2687; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2689 = waySel & _GEN_12211 ? dirty_1_127 : _GEN_2688; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2690 = waySel & _GEN_12213 ? dirty_1_128 : _GEN_2689; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2691 = waySel & _GEN_12215 ? dirty_1_129 : _GEN_2690; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2692 = waySel & _GEN_12217 ? dirty_1_130 : _GEN_2691; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2693 = waySel & _GEN_12219 ? dirty_1_131 : _GEN_2692; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2694 = waySel & _GEN_12221 ? dirty_1_132 : _GEN_2693; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2695 = waySel & _GEN_12223 ? dirty_1_133 : _GEN_2694; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2696 = waySel & _GEN_12225 ? dirty_1_134 : _GEN_2695; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2697 = waySel & _GEN_12227 ? dirty_1_135 : _GEN_2696; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2698 = waySel & _GEN_12229 ? dirty_1_136 : _GEN_2697; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2699 = waySel & _GEN_12231 ? dirty_1_137 : _GEN_2698; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2700 = waySel & _GEN_12233 ? dirty_1_138 : _GEN_2699; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2701 = waySel & _GEN_12235 ? dirty_1_139 : _GEN_2700; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2702 = waySel & _GEN_12237 ? dirty_1_140 : _GEN_2701; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2703 = waySel & _GEN_12239 ? dirty_1_141 : _GEN_2702; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2704 = waySel & _GEN_12241 ? dirty_1_142 : _GEN_2703; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2705 = waySel & _GEN_12243 ? dirty_1_143 : _GEN_2704; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2706 = waySel & _GEN_12245 ? dirty_1_144 : _GEN_2705; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2707 = waySel & _GEN_12247 ? dirty_1_145 : _GEN_2706; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2708 = waySel & _GEN_12249 ? dirty_1_146 : _GEN_2707; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2709 = waySel & _GEN_12251 ? dirty_1_147 : _GEN_2708; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2710 = waySel & _GEN_12253 ? dirty_1_148 : _GEN_2709; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2711 = waySel & _GEN_12255 ? dirty_1_149 : _GEN_2710; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2712 = waySel & _GEN_12257 ? dirty_1_150 : _GEN_2711; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2713 = waySel & _GEN_12259 ? dirty_1_151 : _GEN_2712; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2714 = waySel & _GEN_12261 ? dirty_1_152 : _GEN_2713; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2715 = waySel & _GEN_12263 ? dirty_1_153 : _GEN_2714; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2716 = waySel & _GEN_12265 ? dirty_1_154 : _GEN_2715; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2717 = waySel & _GEN_12267 ? dirty_1_155 : _GEN_2716; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2718 = waySel & _GEN_12269 ? dirty_1_156 : _GEN_2717; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2719 = waySel & _GEN_12271 ? dirty_1_157 : _GEN_2718; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2720 = waySel & _GEN_12273 ? dirty_1_158 : _GEN_2719; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2721 = waySel & _GEN_12275 ? dirty_1_159 : _GEN_2720; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2722 = waySel & _GEN_12277 ? dirty_1_160 : _GEN_2721; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2723 = waySel & _GEN_12279 ? dirty_1_161 : _GEN_2722; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2724 = waySel & _GEN_12281 ? dirty_1_162 : _GEN_2723; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2725 = waySel & _GEN_12283 ? dirty_1_163 : _GEN_2724; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2726 = waySel & _GEN_12285 ? dirty_1_164 : _GEN_2725; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2727 = waySel & _GEN_12287 ? dirty_1_165 : _GEN_2726; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2728 = waySel & _GEN_12289 ? dirty_1_166 : _GEN_2727; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2729 = waySel & _GEN_12291 ? dirty_1_167 : _GEN_2728; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2730 = waySel & _GEN_12293 ? dirty_1_168 : _GEN_2729; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2731 = waySel & _GEN_12295 ? dirty_1_169 : _GEN_2730; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2732 = waySel & _GEN_12297 ? dirty_1_170 : _GEN_2731; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2733 = waySel & _GEN_12299 ? dirty_1_171 : _GEN_2732; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2734 = waySel & _GEN_12301 ? dirty_1_172 : _GEN_2733; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2735 = waySel & _GEN_12303 ? dirty_1_173 : _GEN_2734; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2736 = waySel & _GEN_12305 ? dirty_1_174 : _GEN_2735; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2737 = waySel & _GEN_12307 ? dirty_1_175 : _GEN_2736; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2738 = waySel & _GEN_12309 ? dirty_1_176 : _GEN_2737; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2739 = waySel & _GEN_12311 ? dirty_1_177 : _GEN_2738; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2740 = waySel & _GEN_12313 ? dirty_1_178 : _GEN_2739; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2741 = waySel & _GEN_12315 ? dirty_1_179 : _GEN_2740; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2742 = waySel & _GEN_12317 ? dirty_1_180 : _GEN_2741; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2743 = waySel & _GEN_12319 ? dirty_1_181 : _GEN_2742; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2744 = waySel & _GEN_12321 ? dirty_1_182 : _GEN_2743; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2745 = waySel & _GEN_12323 ? dirty_1_183 : _GEN_2744; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2746 = waySel & _GEN_12325 ? dirty_1_184 : _GEN_2745; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2747 = waySel & _GEN_12327 ? dirty_1_185 : _GEN_2746; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2748 = waySel & _GEN_12329 ? dirty_1_186 : _GEN_2747; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2749 = waySel & _GEN_12331 ? dirty_1_187 : _GEN_2748; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2750 = waySel & _GEN_12333 ? dirty_1_188 : _GEN_2749; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2751 = waySel & _GEN_12335 ? dirty_1_189 : _GEN_2750; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2752 = waySel & _GEN_12337 ? dirty_1_190 : _GEN_2751; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2753 = waySel & _GEN_12339 ? dirty_1_191 : _GEN_2752; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2754 = waySel & _GEN_12341 ? dirty_1_192 : _GEN_2753; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2755 = waySel & _GEN_12343 ? dirty_1_193 : _GEN_2754; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2756 = waySel & _GEN_12345 ? dirty_1_194 : _GEN_2755; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2757 = waySel & _GEN_12347 ? dirty_1_195 : _GEN_2756; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2758 = waySel & _GEN_12349 ? dirty_1_196 : _GEN_2757; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2759 = waySel & _GEN_12351 ? dirty_1_197 : _GEN_2758; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2760 = waySel & _GEN_12353 ? dirty_1_198 : _GEN_2759; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2761 = waySel & _GEN_12355 ? dirty_1_199 : _GEN_2760; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2762 = waySel & _GEN_12357 ? dirty_1_200 : _GEN_2761; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2763 = waySel & _GEN_12359 ? dirty_1_201 : _GEN_2762; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2764 = waySel & _GEN_12361 ? dirty_1_202 : _GEN_2763; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2765 = waySel & _GEN_12363 ? dirty_1_203 : _GEN_2764; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2766 = waySel & _GEN_12365 ? dirty_1_204 : _GEN_2765; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2767 = waySel & _GEN_12367 ? dirty_1_205 : _GEN_2766; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2768 = waySel & _GEN_12369 ? dirty_1_206 : _GEN_2767; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2769 = waySel & _GEN_12371 ? dirty_1_207 : _GEN_2768; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2770 = waySel & _GEN_12373 ? dirty_1_208 : _GEN_2769; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2771 = waySel & _GEN_12375 ? dirty_1_209 : _GEN_2770; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2772 = waySel & _GEN_12377 ? dirty_1_210 : _GEN_2771; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2773 = waySel & _GEN_12379 ? dirty_1_211 : _GEN_2772; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2774 = waySel & _GEN_12381 ? dirty_1_212 : _GEN_2773; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2775 = waySel & _GEN_12383 ? dirty_1_213 : _GEN_2774; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2776 = waySel & _GEN_12385 ? dirty_1_214 : _GEN_2775; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2777 = waySel & _GEN_12387 ? dirty_1_215 : _GEN_2776; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2778 = waySel & _GEN_12389 ? dirty_1_216 : _GEN_2777; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2779 = waySel & _GEN_12391 ? dirty_1_217 : _GEN_2778; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2780 = waySel & _GEN_12393 ? dirty_1_218 : _GEN_2779; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2781 = waySel & _GEN_12395 ? dirty_1_219 : _GEN_2780; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2782 = waySel & _GEN_12397 ? dirty_1_220 : _GEN_2781; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2783 = waySel & _GEN_12399 ? dirty_1_221 : _GEN_2782; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2784 = waySel & _GEN_12401 ? dirty_1_222 : _GEN_2783; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2785 = waySel & _GEN_12403 ? dirty_1_223 : _GEN_2784; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2786 = waySel & _GEN_12405 ? dirty_1_224 : _GEN_2785; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2787 = waySel & _GEN_12407 ? dirty_1_225 : _GEN_2786; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2788 = waySel & _GEN_12409 ? dirty_1_226 : _GEN_2787; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2789 = waySel & _GEN_12411 ? dirty_1_227 : _GEN_2788; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2790 = waySel & _GEN_12413 ? dirty_1_228 : _GEN_2789; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2791 = waySel & _GEN_12415 ? dirty_1_229 : _GEN_2790; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2792 = waySel & _GEN_12417 ? dirty_1_230 : _GEN_2791; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2793 = waySel & _GEN_12419 ? dirty_1_231 : _GEN_2792; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2794 = waySel & _GEN_12421 ? dirty_1_232 : _GEN_2793; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2795 = waySel & _GEN_12423 ? dirty_1_233 : _GEN_2794; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2796 = waySel & _GEN_12425 ? dirty_1_234 : _GEN_2795; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2797 = waySel & _GEN_12427 ? dirty_1_235 : _GEN_2796; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2798 = waySel & _GEN_12429 ? dirty_1_236 : _GEN_2797; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2799 = waySel & _GEN_12431 ? dirty_1_237 : _GEN_2798; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2800 = waySel & _GEN_12433 ? dirty_1_238 : _GEN_2799; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2801 = waySel & _GEN_12435 ? dirty_1_239 : _GEN_2800; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2802 = waySel & _GEN_12437 ? dirty_1_240 : _GEN_2801; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2803 = waySel & _GEN_12439 ? dirty_1_241 : _GEN_2802; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2804 = waySel & _GEN_12441 ? dirty_1_242 : _GEN_2803; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2805 = waySel & _GEN_12443 ? dirty_1_243 : _GEN_2804; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2806 = waySel & _GEN_12445 ? dirty_1_244 : _GEN_2805; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2807 = waySel & _GEN_12447 ? dirty_1_245 : _GEN_2806; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2808 = waySel & _GEN_12449 ? dirty_1_246 : _GEN_2807; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2809 = waySel & _GEN_12451 ? dirty_1_247 : _GEN_2808; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2810 = waySel & _GEN_12453 ? dirty_1_248 : _GEN_2809; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2811 = waySel & _GEN_12455 ? dirty_1_249 : _GEN_2810; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2812 = waySel & _GEN_12457 ? dirty_1_250 : _GEN_2811; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2813 = waySel & _GEN_12459 ? dirty_1_251 : _GEN_2812; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2814 = waySel & _GEN_12461 ? dirty_1_252 : _GEN_2813; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2815 = waySel & _GEN_12463 ? dirty_1_253 : _GEN_2814; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2816 = waySel & _GEN_12465 ? dirty_1_254 : _GEN_2815; // @[Cat.scala 33:{92,92}]
  wire  _GEN_2817 = waySel & _GEN_12467 ? dirty_1_255 : _GEN_2816; // @[Cat.scala 33:{92,92}]
  wire [21:0] _tag_output_T_1 = {_GEN_2817,_GEN_2305}; // @[Cat.scala 33:92]
  wire [21:0] _GEN_2818 = loadTag ? _tag_output_T_1 : 22'h0; // @[dcache.scala 408:30 409:61 98:21]
  wire [20:0] _GEN_2819 = ~waySel ? tag_input[20:0] : 21'h0; // @[dcache.scala 143:25 412:{66,66}]
  wire [20:0] _GEN_2820 = waySel ? tag_input[20:0] : 21'h0; // @[dcache.scala 143:25 412:{66,66}]
  wire  _GEN_2823 = _GEN_13518 & _GEN_12468 ? tag_input[21] : dirty_0_0; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2824 = _GEN_13518 & _GEN_11959 ? tag_input[21] : dirty_0_1; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2825 = _GEN_13518 & _GEN_11961 ? tag_input[21] : dirty_0_2; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2826 = _GEN_13518 & _GEN_11963 ? tag_input[21] : dirty_0_3; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2827 = _GEN_13518 & _GEN_11965 ? tag_input[21] : dirty_0_4; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2828 = _GEN_13518 & _GEN_11967 ? tag_input[21] : dirty_0_5; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2829 = _GEN_13518 & _GEN_11969 ? tag_input[21] : dirty_0_6; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2830 = _GEN_13518 & _GEN_11971 ? tag_input[21] : dirty_0_7; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2831 = _GEN_13518 & _GEN_11973 ? tag_input[21] : dirty_0_8; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2832 = _GEN_13518 & _GEN_11975 ? tag_input[21] : dirty_0_9; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2833 = _GEN_13518 & _GEN_11977 ? tag_input[21] : dirty_0_10; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2834 = _GEN_13518 & _GEN_11979 ? tag_input[21] : dirty_0_11; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2835 = _GEN_13518 & _GEN_11981 ? tag_input[21] : dirty_0_12; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2836 = _GEN_13518 & _GEN_11983 ? tag_input[21] : dirty_0_13; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2837 = _GEN_13518 & _GEN_11985 ? tag_input[21] : dirty_0_14; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2838 = _GEN_13518 & _GEN_11987 ? tag_input[21] : dirty_0_15; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2839 = _GEN_13518 & _GEN_11989 ? tag_input[21] : dirty_0_16; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2840 = _GEN_13518 & _GEN_11991 ? tag_input[21] : dirty_0_17; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2841 = _GEN_13518 & _GEN_11993 ? tag_input[21] : dirty_0_18; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2842 = _GEN_13518 & _GEN_11995 ? tag_input[21] : dirty_0_19; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2843 = _GEN_13518 & _GEN_11997 ? tag_input[21] : dirty_0_20; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2844 = _GEN_13518 & _GEN_11999 ? tag_input[21] : dirty_0_21; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2845 = _GEN_13518 & _GEN_12001 ? tag_input[21] : dirty_0_22; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2846 = _GEN_13518 & _GEN_12003 ? tag_input[21] : dirty_0_23; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2847 = _GEN_13518 & _GEN_12005 ? tag_input[21] : dirty_0_24; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2848 = _GEN_13518 & _GEN_12007 ? tag_input[21] : dirty_0_25; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2849 = _GEN_13518 & _GEN_12009 ? tag_input[21] : dirty_0_26; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2850 = _GEN_13518 & _GEN_12011 ? tag_input[21] : dirty_0_27; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2851 = _GEN_13518 & _GEN_12013 ? tag_input[21] : dirty_0_28; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2852 = _GEN_13518 & _GEN_12015 ? tag_input[21] : dirty_0_29; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2853 = _GEN_13518 & _GEN_12017 ? tag_input[21] : dirty_0_30; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2854 = _GEN_13518 & _GEN_12019 ? tag_input[21] : dirty_0_31; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2855 = _GEN_13518 & _GEN_12021 ? tag_input[21] : dirty_0_32; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2856 = _GEN_13518 & _GEN_12023 ? tag_input[21] : dirty_0_33; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2857 = _GEN_13518 & _GEN_12025 ? tag_input[21] : dirty_0_34; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2858 = _GEN_13518 & _GEN_12027 ? tag_input[21] : dirty_0_35; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2859 = _GEN_13518 & _GEN_12029 ? tag_input[21] : dirty_0_36; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2860 = _GEN_13518 & _GEN_12031 ? tag_input[21] : dirty_0_37; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2861 = _GEN_13518 & _GEN_12033 ? tag_input[21] : dirty_0_38; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2862 = _GEN_13518 & _GEN_12035 ? tag_input[21] : dirty_0_39; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2863 = _GEN_13518 & _GEN_12037 ? tag_input[21] : dirty_0_40; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2864 = _GEN_13518 & _GEN_12039 ? tag_input[21] : dirty_0_41; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2865 = _GEN_13518 & _GEN_12041 ? tag_input[21] : dirty_0_42; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2866 = _GEN_13518 & _GEN_12043 ? tag_input[21] : dirty_0_43; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2867 = _GEN_13518 & _GEN_12045 ? tag_input[21] : dirty_0_44; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2868 = _GEN_13518 & _GEN_12047 ? tag_input[21] : dirty_0_45; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2869 = _GEN_13518 & _GEN_12049 ? tag_input[21] : dirty_0_46; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2870 = _GEN_13518 & _GEN_12051 ? tag_input[21] : dirty_0_47; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2871 = _GEN_13518 & _GEN_12053 ? tag_input[21] : dirty_0_48; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2872 = _GEN_13518 & _GEN_12055 ? tag_input[21] : dirty_0_49; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2873 = _GEN_13518 & _GEN_12057 ? tag_input[21] : dirty_0_50; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2874 = _GEN_13518 & _GEN_12059 ? tag_input[21] : dirty_0_51; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2875 = _GEN_13518 & _GEN_12061 ? tag_input[21] : dirty_0_52; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2876 = _GEN_13518 & _GEN_12063 ? tag_input[21] : dirty_0_53; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2877 = _GEN_13518 & _GEN_12065 ? tag_input[21] : dirty_0_54; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2878 = _GEN_13518 & _GEN_12067 ? tag_input[21] : dirty_0_55; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2879 = _GEN_13518 & _GEN_12069 ? tag_input[21] : dirty_0_56; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2880 = _GEN_13518 & _GEN_12071 ? tag_input[21] : dirty_0_57; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2881 = _GEN_13518 & _GEN_12073 ? tag_input[21] : dirty_0_58; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2882 = _GEN_13518 & _GEN_12075 ? tag_input[21] : dirty_0_59; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2883 = _GEN_13518 & _GEN_12077 ? tag_input[21] : dirty_0_60; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2884 = _GEN_13518 & _GEN_12079 ? tag_input[21] : dirty_0_61; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2885 = _GEN_13518 & _GEN_12081 ? tag_input[21] : dirty_0_62; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2886 = _GEN_13518 & _GEN_12083 ? tag_input[21] : dirty_0_63; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2887 = _GEN_13518 & _GEN_12085 ? tag_input[21] : dirty_0_64; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2888 = _GEN_13518 & _GEN_12087 ? tag_input[21] : dirty_0_65; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2889 = _GEN_13518 & _GEN_12089 ? tag_input[21] : dirty_0_66; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2890 = _GEN_13518 & _GEN_12091 ? tag_input[21] : dirty_0_67; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2891 = _GEN_13518 & _GEN_12093 ? tag_input[21] : dirty_0_68; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2892 = _GEN_13518 & _GEN_12095 ? tag_input[21] : dirty_0_69; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2893 = _GEN_13518 & _GEN_12097 ? tag_input[21] : dirty_0_70; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2894 = _GEN_13518 & _GEN_12099 ? tag_input[21] : dirty_0_71; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2895 = _GEN_13518 & _GEN_12101 ? tag_input[21] : dirty_0_72; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2896 = _GEN_13518 & _GEN_12103 ? tag_input[21] : dirty_0_73; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2897 = _GEN_13518 & _GEN_12105 ? tag_input[21] : dirty_0_74; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2898 = _GEN_13518 & _GEN_12107 ? tag_input[21] : dirty_0_75; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2899 = _GEN_13518 & _GEN_12109 ? tag_input[21] : dirty_0_76; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2900 = _GEN_13518 & _GEN_12111 ? tag_input[21] : dirty_0_77; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2901 = _GEN_13518 & _GEN_12113 ? tag_input[21] : dirty_0_78; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2902 = _GEN_13518 & _GEN_12115 ? tag_input[21] : dirty_0_79; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2903 = _GEN_13518 & _GEN_12117 ? tag_input[21] : dirty_0_80; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2904 = _GEN_13518 & _GEN_12119 ? tag_input[21] : dirty_0_81; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2905 = _GEN_13518 & _GEN_12121 ? tag_input[21] : dirty_0_82; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2906 = _GEN_13518 & _GEN_12123 ? tag_input[21] : dirty_0_83; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2907 = _GEN_13518 & _GEN_12125 ? tag_input[21] : dirty_0_84; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2908 = _GEN_13518 & _GEN_12127 ? tag_input[21] : dirty_0_85; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2909 = _GEN_13518 & _GEN_12129 ? tag_input[21] : dirty_0_86; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2910 = _GEN_13518 & _GEN_12131 ? tag_input[21] : dirty_0_87; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2911 = _GEN_13518 & _GEN_12133 ? tag_input[21] : dirty_0_88; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2912 = _GEN_13518 & _GEN_12135 ? tag_input[21] : dirty_0_89; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2913 = _GEN_13518 & _GEN_12137 ? tag_input[21] : dirty_0_90; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2914 = _GEN_13518 & _GEN_12139 ? tag_input[21] : dirty_0_91; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2915 = _GEN_13518 & _GEN_12141 ? tag_input[21] : dirty_0_92; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2916 = _GEN_13518 & _GEN_12143 ? tag_input[21] : dirty_0_93; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2917 = _GEN_13518 & _GEN_12145 ? tag_input[21] : dirty_0_94; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2918 = _GEN_13518 & _GEN_12147 ? tag_input[21] : dirty_0_95; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2919 = _GEN_13518 & _GEN_12149 ? tag_input[21] : dirty_0_96; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2920 = _GEN_13518 & _GEN_12151 ? tag_input[21] : dirty_0_97; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2921 = _GEN_13518 & _GEN_12153 ? tag_input[21] : dirty_0_98; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2922 = _GEN_13518 & _GEN_12155 ? tag_input[21] : dirty_0_99; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2923 = _GEN_13518 & _GEN_12157 ? tag_input[21] : dirty_0_100; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2924 = _GEN_13518 & _GEN_12159 ? tag_input[21] : dirty_0_101; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2925 = _GEN_13518 & _GEN_12161 ? tag_input[21] : dirty_0_102; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2926 = _GEN_13518 & _GEN_12163 ? tag_input[21] : dirty_0_103; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2927 = _GEN_13518 & _GEN_12165 ? tag_input[21] : dirty_0_104; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2928 = _GEN_13518 & _GEN_12167 ? tag_input[21] : dirty_0_105; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2929 = _GEN_13518 & _GEN_12169 ? tag_input[21] : dirty_0_106; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2930 = _GEN_13518 & _GEN_12171 ? tag_input[21] : dirty_0_107; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2931 = _GEN_13518 & _GEN_12173 ? tag_input[21] : dirty_0_108; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2932 = _GEN_13518 & _GEN_12175 ? tag_input[21] : dirty_0_109; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2933 = _GEN_13518 & _GEN_12177 ? tag_input[21] : dirty_0_110; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2934 = _GEN_13518 & _GEN_12179 ? tag_input[21] : dirty_0_111; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2935 = _GEN_13518 & _GEN_12181 ? tag_input[21] : dirty_0_112; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2936 = _GEN_13518 & _GEN_12183 ? tag_input[21] : dirty_0_113; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2937 = _GEN_13518 & _GEN_12185 ? tag_input[21] : dirty_0_114; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2938 = _GEN_13518 & _GEN_12187 ? tag_input[21] : dirty_0_115; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2939 = _GEN_13518 & _GEN_12189 ? tag_input[21] : dirty_0_116; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2940 = _GEN_13518 & _GEN_12191 ? tag_input[21] : dirty_0_117; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2941 = _GEN_13518 & _GEN_12193 ? tag_input[21] : dirty_0_118; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2942 = _GEN_13518 & _GEN_12195 ? tag_input[21] : dirty_0_119; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2943 = _GEN_13518 & _GEN_12197 ? tag_input[21] : dirty_0_120; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2944 = _GEN_13518 & _GEN_12199 ? tag_input[21] : dirty_0_121; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2945 = _GEN_13518 & _GEN_12201 ? tag_input[21] : dirty_0_122; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2946 = _GEN_13518 & _GEN_12203 ? tag_input[21] : dirty_0_123; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2947 = _GEN_13518 & _GEN_12205 ? tag_input[21] : dirty_0_124; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2948 = _GEN_13518 & _GEN_12207 ? tag_input[21] : dirty_0_125; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2949 = _GEN_13518 & _GEN_12209 ? tag_input[21] : dirty_0_126; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2950 = _GEN_13518 & _GEN_12211 ? tag_input[21] : dirty_0_127; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2951 = _GEN_13518 & _GEN_12213 ? tag_input[21] : dirty_0_128; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2952 = _GEN_13518 & _GEN_12215 ? tag_input[21] : dirty_0_129; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2953 = _GEN_13518 & _GEN_12217 ? tag_input[21] : dirty_0_130; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2954 = _GEN_13518 & _GEN_12219 ? tag_input[21] : dirty_0_131; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2955 = _GEN_13518 & _GEN_12221 ? tag_input[21] : dirty_0_132; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2956 = _GEN_13518 & _GEN_12223 ? tag_input[21] : dirty_0_133; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2957 = _GEN_13518 & _GEN_12225 ? tag_input[21] : dirty_0_134; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2958 = _GEN_13518 & _GEN_12227 ? tag_input[21] : dirty_0_135; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2959 = _GEN_13518 & _GEN_12229 ? tag_input[21] : dirty_0_136; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2960 = _GEN_13518 & _GEN_12231 ? tag_input[21] : dirty_0_137; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2961 = _GEN_13518 & _GEN_12233 ? tag_input[21] : dirty_0_138; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2962 = _GEN_13518 & _GEN_12235 ? tag_input[21] : dirty_0_139; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2963 = _GEN_13518 & _GEN_12237 ? tag_input[21] : dirty_0_140; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2964 = _GEN_13518 & _GEN_12239 ? tag_input[21] : dirty_0_141; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2965 = _GEN_13518 & _GEN_12241 ? tag_input[21] : dirty_0_142; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2966 = _GEN_13518 & _GEN_12243 ? tag_input[21] : dirty_0_143; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2967 = _GEN_13518 & _GEN_12245 ? tag_input[21] : dirty_0_144; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2968 = _GEN_13518 & _GEN_12247 ? tag_input[21] : dirty_0_145; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2969 = _GEN_13518 & _GEN_12249 ? tag_input[21] : dirty_0_146; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2970 = _GEN_13518 & _GEN_12251 ? tag_input[21] : dirty_0_147; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2971 = _GEN_13518 & _GEN_12253 ? tag_input[21] : dirty_0_148; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2972 = _GEN_13518 & _GEN_12255 ? tag_input[21] : dirty_0_149; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2973 = _GEN_13518 & _GEN_12257 ? tag_input[21] : dirty_0_150; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2974 = _GEN_13518 & _GEN_12259 ? tag_input[21] : dirty_0_151; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2975 = _GEN_13518 & _GEN_12261 ? tag_input[21] : dirty_0_152; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2976 = _GEN_13518 & _GEN_12263 ? tag_input[21] : dirty_0_153; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2977 = _GEN_13518 & _GEN_12265 ? tag_input[21] : dirty_0_154; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2978 = _GEN_13518 & _GEN_12267 ? tag_input[21] : dirty_0_155; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2979 = _GEN_13518 & _GEN_12269 ? tag_input[21] : dirty_0_156; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2980 = _GEN_13518 & _GEN_12271 ? tag_input[21] : dirty_0_157; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2981 = _GEN_13518 & _GEN_12273 ? tag_input[21] : dirty_0_158; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2982 = _GEN_13518 & _GEN_12275 ? tag_input[21] : dirty_0_159; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2983 = _GEN_13518 & _GEN_12277 ? tag_input[21] : dirty_0_160; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2984 = _GEN_13518 & _GEN_12279 ? tag_input[21] : dirty_0_161; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2985 = _GEN_13518 & _GEN_12281 ? tag_input[21] : dirty_0_162; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2986 = _GEN_13518 & _GEN_12283 ? tag_input[21] : dirty_0_163; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2987 = _GEN_13518 & _GEN_12285 ? tag_input[21] : dirty_0_164; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2988 = _GEN_13518 & _GEN_12287 ? tag_input[21] : dirty_0_165; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2989 = _GEN_13518 & _GEN_12289 ? tag_input[21] : dirty_0_166; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2990 = _GEN_13518 & _GEN_12291 ? tag_input[21] : dirty_0_167; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2991 = _GEN_13518 & _GEN_12293 ? tag_input[21] : dirty_0_168; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2992 = _GEN_13518 & _GEN_12295 ? tag_input[21] : dirty_0_169; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2993 = _GEN_13518 & _GEN_12297 ? tag_input[21] : dirty_0_170; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2994 = _GEN_13518 & _GEN_12299 ? tag_input[21] : dirty_0_171; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2995 = _GEN_13518 & _GEN_12301 ? tag_input[21] : dirty_0_172; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2996 = _GEN_13518 & _GEN_12303 ? tag_input[21] : dirty_0_173; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2997 = _GEN_13518 & _GEN_12305 ? tag_input[21] : dirty_0_174; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2998 = _GEN_13518 & _GEN_12307 ? tag_input[21] : dirty_0_175; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_2999 = _GEN_13518 & _GEN_12309 ? tag_input[21] : dirty_0_176; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3000 = _GEN_13518 & _GEN_12311 ? tag_input[21] : dirty_0_177; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3001 = _GEN_13518 & _GEN_12313 ? tag_input[21] : dirty_0_178; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3002 = _GEN_13518 & _GEN_12315 ? tag_input[21] : dirty_0_179; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3003 = _GEN_13518 & _GEN_12317 ? tag_input[21] : dirty_0_180; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3004 = _GEN_13518 & _GEN_12319 ? tag_input[21] : dirty_0_181; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3005 = _GEN_13518 & _GEN_12321 ? tag_input[21] : dirty_0_182; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3006 = _GEN_13518 & _GEN_12323 ? tag_input[21] : dirty_0_183; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3007 = _GEN_13518 & _GEN_12325 ? tag_input[21] : dirty_0_184; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3008 = _GEN_13518 & _GEN_12327 ? tag_input[21] : dirty_0_185; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3009 = _GEN_13518 & _GEN_12329 ? tag_input[21] : dirty_0_186; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3010 = _GEN_13518 & _GEN_12331 ? tag_input[21] : dirty_0_187; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3011 = _GEN_13518 & _GEN_12333 ? tag_input[21] : dirty_0_188; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3012 = _GEN_13518 & _GEN_12335 ? tag_input[21] : dirty_0_189; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3013 = _GEN_13518 & _GEN_12337 ? tag_input[21] : dirty_0_190; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3014 = _GEN_13518 & _GEN_12339 ? tag_input[21] : dirty_0_191; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3015 = _GEN_13518 & _GEN_12341 ? tag_input[21] : dirty_0_192; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3016 = _GEN_13518 & _GEN_12343 ? tag_input[21] : dirty_0_193; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3017 = _GEN_13518 & _GEN_12345 ? tag_input[21] : dirty_0_194; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3018 = _GEN_13518 & _GEN_12347 ? tag_input[21] : dirty_0_195; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3019 = _GEN_13518 & _GEN_12349 ? tag_input[21] : dirty_0_196; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3020 = _GEN_13518 & _GEN_12351 ? tag_input[21] : dirty_0_197; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3021 = _GEN_13518 & _GEN_12353 ? tag_input[21] : dirty_0_198; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3022 = _GEN_13518 & _GEN_12355 ? tag_input[21] : dirty_0_199; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3023 = _GEN_13518 & _GEN_12357 ? tag_input[21] : dirty_0_200; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3024 = _GEN_13518 & _GEN_12359 ? tag_input[21] : dirty_0_201; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3025 = _GEN_13518 & _GEN_12361 ? tag_input[21] : dirty_0_202; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3026 = _GEN_13518 & _GEN_12363 ? tag_input[21] : dirty_0_203; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3027 = _GEN_13518 & _GEN_12365 ? tag_input[21] : dirty_0_204; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3028 = _GEN_13518 & _GEN_12367 ? tag_input[21] : dirty_0_205; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3029 = _GEN_13518 & _GEN_12369 ? tag_input[21] : dirty_0_206; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3030 = _GEN_13518 & _GEN_12371 ? tag_input[21] : dirty_0_207; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3031 = _GEN_13518 & _GEN_12373 ? tag_input[21] : dirty_0_208; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3032 = _GEN_13518 & _GEN_12375 ? tag_input[21] : dirty_0_209; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3033 = _GEN_13518 & _GEN_12377 ? tag_input[21] : dirty_0_210; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3034 = _GEN_13518 & _GEN_12379 ? tag_input[21] : dirty_0_211; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3035 = _GEN_13518 & _GEN_12381 ? tag_input[21] : dirty_0_212; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3036 = _GEN_13518 & _GEN_12383 ? tag_input[21] : dirty_0_213; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3037 = _GEN_13518 & _GEN_12385 ? tag_input[21] : dirty_0_214; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3038 = _GEN_13518 & _GEN_12387 ? tag_input[21] : dirty_0_215; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3039 = _GEN_13518 & _GEN_12389 ? tag_input[21] : dirty_0_216; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3040 = _GEN_13518 & _GEN_12391 ? tag_input[21] : dirty_0_217; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3041 = _GEN_13518 & _GEN_12393 ? tag_input[21] : dirty_0_218; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3042 = _GEN_13518 & _GEN_12395 ? tag_input[21] : dirty_0_219; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3043 = _GEN_13518 & _GEN_12397 ? tag_input[21] : dirty_0_220; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3044 = _GEN_13518 & _GEN_12399 ? tag_input[21] : dirty_0_221; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3045 = _GEN_13518 & _GEN_12401 ? tag_input[21] : dirty_0_222; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3046 = _GEN_13518 & _GEN_12403 ? tag_input[21] : dirty_0_223; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3047 = _GEN_13518 & _GEN_12405 ? tag_input[21] : dirty_0_224; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3048 = _GEN_13518 & _GEN_12407 ? tag_input[21] : dirty_0_225; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3049 = _GEN_13518 & _GEN_12409 ? tag_input[21] : dirty_0_226; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3050 = _GEN_13518 & _GEN_12411 ? tag_input[21] : dirty_0_227; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3051 = _GEN_13518 & _GEN_12413 ? tag_input[21] : dirty_0_228; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3052 = _GEN_13518 & _GEN_12415 ? tag_input[21] : dirty_0_229; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3053 = _GEN_13518 & _GEN_12417 ? tag_input[21] : dirty_0_230; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3054 = _GEN_13518 & _GEN_12419 ? tag_input[21] : dirty_0_231; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3055 = _GEN_13518 & _GEN_12421 ? tag_input[21] : dirty_0_232; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3056 = _GEN_13518 & _GEN_12423 ? tag_input[21] : dirty_0_233; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3057 = _GEN_13518 & _GEN_12425 ? tag_input[21] : dirty_0_234; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3058 = _GEN_13518 & _GEN_12427 ? tag_input[21] : dirty_0_235; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3059 = _GEN_13518 & _GEN_12429 ? tag_input[21] : dirty_0_236; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3060 = _GEN_13518 & _GEN_12431 ? tag_input[21] : dirty_0_237; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3061 = _GEN_13518 & _GEN_12433 ? tag_input[21] : dirty_0_238; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3062 = _GEN_13518 & _GEN_12435 ? tag_input[21] : dirty_0_239; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3063 = _GEN_13518 & _GEN_12437 ? tag_input[21] : dirty_0_240; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3064 = _GEN_13518 & _GEN_12439 ? tag_input[21] : dirty_0_241; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3065 = _GEN_13518 & _GEN_12441 ? tag_input[21] : dirty_0_242; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3066 = _GEN_13518 & _GEN_12443 ? tag_input[21] : dirty_0_243; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3067 = _GEN_13518 & _GEN_12445 ? tag_input[21] : dirty_0_244; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3068 = _GEN_13518 & _GEN_12447 ? tag_input[21] : dirty_0_245; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3069 = _GEN_13518 & _GEN_12449 ? tag_input[21] : dirty_0_246; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3070 = _GEN_13518 & _GEN_12451 ? tag_input[21] : dirty_0_247; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3071 = _GEN_13518 & _GEN_12453 ? tag_input[21] : dirty_0_248; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3072 = _GEN_13518 & _GEN_12455 ? tag_input[21] : dirty_0_249; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3073 = _GEN_13518 & _GEN_12457 ? tag_input[21] : dirty_0_250; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3074 = _GEN_13518 & _GEN_12459 ? tag_input[21] : dirty_0_251; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3075 = _GEN_13518 & _GEN_12461 ? tag_input[21] : dirty_0_252; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3076 = _GEN_13518 & _GEN_12463 ? tag_input[21] : dirty_0_253; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3077 = _GEN_13518 & _GEN_12465 ? tag_input[21] : dirty_0_254; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3078 = _GEN_13518 & _GEN_12467 ? tag_input[21] : dirty_0_255; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3079 = waySel & _GEN_12468 ? tag_input[21] : dirty_1_0; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3080 = waySel & _GEN_11959 ? tag_input[21] : dirty_1_1; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3081 = waySel & _GEN_11961 ? tag_input[21] : dirty_1_2; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3082 = waySel & _GEN_11963 ? tag_input[21] : dirty_1_3; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3083 = waySel & _GEN_11965 ? tag_input[21] : dirty_1_4; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3084 = waySel & _GEN_11967 ? tag_input[21] : dirty_1_5; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3085 = waySel & _GEN_11969 ? tag_input[21] : dirty_1_6; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3086 = waySel & _GEN_11971 ? tag_input[21] : dirty_1_7; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3087 = waySel & _GEN_11973 ? tag_input[21] : dirty_1_8; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3088 = waySel & _GEN_11975 ? tag_input[21] : dirty_1_9; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3089 = waySel & _GEN_11977 ? tag_input[21] : dirty_1_10; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3090 = waySel & _GEN_11979 ? tag_input[21] : dirty_1_11; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3091 = waySel & _GEN_11981 ? tag_input[21] : dirty_1_12; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3092 = waySel & _GEN_11983 ? tag_input[21] : dirty_1_13; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3093 = waySel & _GEN_11985 ? tag_input[21] : dirty_1_14; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3094 = waySel & _GEN_11987 ? tag_input[21] : dirty_1_15; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3095 = waySel & _GEN_11989 ? tag_input[21] : dirty_1_16; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3096 = waySel & _GEN_11991 ? tag_input[21] : dirty_1_17; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3097 = waySel & _GEN_11993 ? tag_input[21] : dirty_1_18; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3098 = waySel & _GEN_11995 ? tag_input[21] : dirty_1_19; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3099 = waySel & _GEN_11997 ? tag_input[21] : dirty_1_20; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3100 = waySel & _GEN_11999 ? tag_input[21] : dirty_1_21; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3101 = waySel & _GEN_12001 ? tag_input[21] : dirty_1_22; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3102 = waySel & _GEN_12003 ? tag_input[21] : dirty_1_23; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3103 = waySel & _GEN_12005 ? tag_input[21] : dirty_1_24; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3104 = waySel & _GEN_12007 ? tag_input[21] : dirty_1_25; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3105 = waySel & _GEN_12009 ? tag_input[21] : dirty_1_26; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3106 = waySel & _GEN_12011 ? tag_input[21] : dirty_1_27; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3107 = waySel & _GEN_12013 ? tag_input[21] : dirty_1_28; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3108 = waySel & _GEN_12015 ? tag_input[21] : dirty_1_29; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3109 = waySel & _GEN_12017 ? tag_input[21] : dirty_1_30; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3110 = waySel & _GEN_12019 ? tag_input[21] : dirty_1_31; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3111 = waySel & _GEN_12021 ? tag_input[21] : dirty_1_32; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3112 = waySel & _GEN_12023 ? tag_input[21] : dirty_1_33; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3113 = waySel & _GEN_12025 ? tag_input[21] : dirty_1_34; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3114 = waySel & _GEN_12027 ? tag_input[21] : dirty_1_35; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3115 = waySel & _GEN_12029 ? tag_input[21] : dirty_1_36; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3116 = waySel & _GEN_12031 ? tag_input[21] : dirty_1_37; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3117 = waySel & _GEN_12033 ? tag_input[21] : dirty_1_38; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3118 = waySel & _GEN_12035 ? tag_input[21] : dirty_1_39; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3119 = waySel & _GEN_12037 ? tag_input[21] : dirty_1_40; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3120 = waySel & _GEN_12039 ? tag_input[21] : dirty_1_41; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3121 = waySel & _GEN_12041 ? tag_input[21] : dirty_1_42; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3122 = waySel & _GEN_12043 ? tag_input[21] : dirty_1_43; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3123 = waySel & _GEN_12045 ? tag_input[21] : dirty_1_44; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3124 = waySel & _GEN_12047 ? tag_input[21] : dirty_1_45; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3125 = waySel & _GEN_12049 ? tag_input[21] : dirty_1_46; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3126 = waySel & _GEN_12051 ? tag_input[21] : dirty_1_47; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3127 = waySel & _GEN_12053 ? tag_input[21] : dirty_1_48; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3128 = waySel & _GEN_12055 ? tag_input[21] : dirty_1_49; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3129 = waySel & _GEN_12057 ? tag_input[21] : dirty_1_50; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3130 = waySel & _GEN_12059 ? tag_input[21] : dirty_1_51; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3131 = waySel & _GEN_12061 ? tag_input[21] : dirty_1_52; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3132 = waySel & _GEN_12063 ? tag_input[21] : dirty_1_53; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3133 = waySel & _GEN_12065 ? tag_input[21] : dirty_1_54; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3134 = waySel & _GEN_12067 ? tag_input[21] : dirty_1_55; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3135 = waySel & _GEN_12069 ? tag_input[21] : dirty_1_56; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3136 = waySel & _GEN_12071 ? tag_input[21] : dirty_1_57; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3137 = waySel & _GEN_12073 ? tag_input[21] : dirty_1_58; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3138 = waySel & _GEN_12075 ? tag_input[21] : dirty_1_59; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3139 = waySel & _GEN_12077 ? tag_input[21] : dirty_1_60; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3140 = waySel & _GEN_12079 ? tag_input[21] : dirty_1_61; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3141 = waySel & _GEN_12081 ? tag_input[21] : dirty_1_62; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3142 = waySel & _GEN_12083 ? tag_input[21] : dirty_1_63; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3143 = waySel & _GEN_12085 ? tag_input[21] : dirty_1_64; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3144 = waySel & _GEN_12087 ? tag_input[21] : dirty_1_65; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3145 = waySel & _GEN_12089 ? tag_input[21] : dirty_1_66; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3146 = waySel & _GEN_12091 ? tag_input[21] : dirty_1_67; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3147 = waySel & _GEN_12093 ? tag_input[21] : dirty_1_68; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3148 = waySel & _GEN_12095 ? tag_input[21] : dirty_1_69; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3149 = waySel & _GEN_12097 ? tag_input[21] : dirty_1_70; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3150 = waySel & _GEN_12099 ? tag_input[21] : dirty_1_71; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3151 = waySel & _GEN_12101 ? tag_input[21] : dirty_1_72; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3152 = waySel & _GEN_12103 ? tag_input[21] : dirty_1_73; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3153 = waySel & _GEN_12105 ? tag_input[21] : dirty_1_74; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3154 = waySel & _GEN_12107 ? tag_input[21] : dirty_1_75; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3155 = waySel & _GEN_12109 ? tag_input[21] : dirty_1_76; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3156 = waySel & _GEN_12111 ? tag_input[21] : dirty_1_77; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3157 = waySel & _GEN_12113 ? tag_input[21] : dirty_1_78; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3158 = waySel & _GEN_12115 ? tag_input[21] : dirty_1_79; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3159 = waySel & _GEN_12117 ? tag_input[21] : dirty_1_80; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3160 = waySel & _GEN_12119 ? tag_input[21] : dirty_1_81; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3161 = waySel & _GEN_12121 ? tag_input[21] : dirty_1_82; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3162 = waySel & _GEN_12123 ? tag_input[21] : dirty_1_83; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3163 = waySel & _GEN_12125 ? tag_input[21] : dirty_1_84; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3164 = waySel & _GEN_12127 ? tag_input[21] : dirty_1_85; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3165 = waySel & _GEN_12129 ? tag_input[21] : dirty_1_86; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3166 = waySel & _GEN_12131 ? tag_input[21] : dirty_1_87; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3167 = waySel & _GEN_12133 ? tag_input[21] : dirty_1_88; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3168 = waySel & _GEN_12135 ? tag_input[21] : dirty_1_89; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3169 = waySel & _GEN_12137 ? tag_input[21] : dirty_1_90; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3170 = waySel & _GEN_12139 ? tag_input[21] : dirty_1_91; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3171 = waySel & _GEN_12141 ? tag_input[21] : dirty_1_92; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3172 = waySel & _GEN_12143 ? tag_input[21] : dirty_1_93; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3173 = waySel & _GEN_12145 ? tag_input[21] : dirty_1_94; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3174 = waySel & _GEN_12147 ? tag_input[21] : dirty_1_95; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3175 = waySel & _GEN_12149 ? tag_input[21] : dirty_1_96; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3176 = waySel & _GEN_12151 ? tag_input[21] : dirty_1_97; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3177 = waySel & _GEN_12153 ? tag_input[21] : dirty_1_98; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3178 = waySel & _GEN_12155 ? tag_input[21] : dirty_1_99; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3179 = waySel & _GEN_12157 ? tag_input[21] : dirty_1_100; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3180 = waySel & _GEN_12159 ? tag_input[21] : dirty_1_101; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3181 = waySel & _GEN_12161 ? tag_input[21] : dirty_1_102; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3182 = waySel & _GEN_12163 ? tag_input[21] : dirty_1_103; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3183 = waySel & _GEN_12165 ? tag_input[21] : dirty_1_104; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3184 = waySel & _GEN_12167 ? tag_input[21] : dirty_1_105; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3185 = waySel & _GEN_12169 ? tag_input[21] : dirty_1_106; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3186 = waySel & _GEN_12171 ? tag_input[21] : dirty_1_107; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3187 = waySel & _GEN_12173 ? tag_input[21] : dirty_1_108; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3188 = waySel & _GEN_12175 ? tag_input[21] : dirty_1_109; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3189 = waySel & _GEN_12177 ? tag_input[21] : dirty_1_110; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3190 = waySel & _GEN_12179 ? tag_input[21] : dirty_1_111; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3191 = waySel & _GEN_12181 ? tag_input[21] : dirty_1_112; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3192 = waySel & _GEN_12183 ? tag_input[21] : dirty_1_113; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3193 = waySel & _GEN_12185 ? tag_input[21] : dirty_1_114; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3194 = waySel & _GEN_12187 ? tag_input[21] : dirty_1_115; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3195 = waySel & _GEN_12189 ? tag_input[21] : dirty_1_116; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3196 = waySel & _GEN_12191 ? tag_input[21] : dirty_1_117; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3197 = waySel & _GEN_12193 ? tag_input[21] : dirty_1_118; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3198 = waySel & _GEN_12195 ? tag_input[21] : dirty_1_119; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3199 = waySel & _GEN_12197 ? tag_input[21] : dirty_1_120; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3200 = waySel & _GEN_12199 ? tag_input[21] : dirty_1_121; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3201 = waySel & _GEN_12201 ? tag_input[21] : dirty_1_122; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3202 = waySel & _GEN_12203 ? tag_input[21] : dirty_1_123; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3203 = waySel & _GEN_12205 ? tag_input[21] : dirty_1_124; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3204 = waySel & _GEN_12207 ? tag_input[21] : dirty_1_125; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3205 = waySel & _GEN_12209 ? tag_input[21] : dirty_1_126; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3206 = waySel & _GEN_12211 ? tag_input[21] : dirty_1_127; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3207 = waySel & _GEN_12213 ? tag_input[21] : dirty_1_128; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3208 = waySel & _GEN_12215 ? tag_input[21] : dirty_1_129; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3209 = waySel & _GEN_12217 ? tag_input[21] : dirty_1_130; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3210 = waySel & _GEN_12219 ? tag_input[21] : dirty_1_131; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3211 = waySel & _GEN_12221 ? tag_input[21] : dirty_1_132; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3212 = waySel & _GEN_12223 ? tag_input[21] : dirty_1_133; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3213 = waySel & _GEN_12225 ? tag_input[21] : dirty_1_134; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3214 = waySel & _GEN_12227 ? tag_input[21] : dirty_1_135; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3215 = waySel & _GEN_12229 ? tag_input[21] : dirty_1_136; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3216 = waySel & _GEN_12231 ? tag_input[21] : dirty_1_137; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3217 = waySel & _GEN_12233 ? tag_input[21] : dirty_1_138; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3218 = waySel & _GEN_12235 ? tag_input[21] : dirty_1_139; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3219 = waySel & _GEN_12237 ? tag_input[21] : dirty_1_140; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3220 = waySel & _GEN_12239 ? tag_input[21] : dirty_1_141; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3221 = waySel & _GEN_12241 ? tag_input[21] : dirty_1_142; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3222 = waySel & _GEN_12243 ? tag_input[21] : dirty_1_143; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3223 = waySel & _GEN_12245 ? tag_input[21] : dirty_1_144; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3224 = waySel & _GEN_12247 ? tag_input[21] : dirty_1_145; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3225 = waySel & _GEN_12249 ? tag_input[21] : dirty_1_146; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3226 = waySel & _GEN_12251 ? tag_input[21] : dirty_1_147; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3227 = waySel & _GEN_12253 ? tag_input[21] : dirty_1_148; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3228 = waySel & _GEN_12255 ? tag_input[21] : dirty_1_149; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3229 = waySel & _GEN_12257 ? tag_input[21] : dirty_1_150; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3230 = waySel & _GEN_12259 ? tag_input[21] : dirty_1_151; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3231 = waySel & _GEN_12261 ? tag_input[21] : dirty_1_152; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3232 = waySel & _GEN_12263 ? tag_input[21] : dirty_1_153; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3233 = waySel & _GEN_12265 ? tag_input[21] : dirty_1_154; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3234 = waySel & _GEN_12267 ? tag_input[21] : dirty_1_155; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3235 = waySel & _GEN_12269 ? tag_input[21] : dirty_1_156; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3236 = waySel & _GEN_12271 ? tag_input[21] : dirty_1_157; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3237 = waySel & _GEN_12273 ? tag_input[21] : dirty_1_158; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3238 = waySel & _GEN_12275 ? tag_input[21] : dirty_1_159; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3239 = waySel & _GEN_12277 ? tag_input[21] : dirty_1_160; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3240 = waySel & _GEN_12279 ? tag_input[21] : dirty_1_161; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3241 = waySel & _GEN_12281 ? tag_input[21] : dirty_1_162; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3242 = waySel & _GEN_12283 ? tag_input[21] : dirty_1_163; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3243 = waySel & _GEN_12285 ? tag_input[21] : dirty_1_164; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3244 = waySel & _GEN_12287 ? tag_input[21] : dirty_1_165; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3245 = waySel & _GEN_12289 ? tag_input[21] : dirty_1_166; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3246 = waySel & _GEN_12291 ? tag_input[21] : dirty_1_167; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3247 = waySel & _GEN_12293 ? tag_input[21] : dirty_1_168; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3248 = waySel & _GEN_12295 ? tag_input[21] : dirty_1_169; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3249 = waySel & _GEN_12297 ? tag_input[21] : dirty_1_170; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3250 = waySel & _GEN_12299 ? tag_input[21] : dirty_1_171; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3251 = waySel & _GEN_12301 ? tag_input[21] : dirty_1_172; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3252 = waySel & _GEN_12303 ? tag_input[21] : dirty_1_173; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3253 = waySel & _GEN_12305 ? tag_input[21] : dirty_1_174; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3254 = waySel & _GEN_12307 ? tag_input[21] : dirty_1_175; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3255 = waySel & _GEN_12309 ? tag_input[21] : dirty_1_176; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3256 = waySel & _GEN_12311 ? tag_input[21] : dirty_1_177; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3257 = waySel & _GEN_12313 ? tag_input[21] : dirty_1_178; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3258 = waySel & _GEN_12315 ? tag_input[21] : dirty_1_179; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3259 = waySel & _GEN_12317 ? tag_input[21] : dirty_1_180; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3260 = waySel & _GEN_12319 ? tag_input[21] : dirty_1_181; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3261 = waySel & _GEN_12321 ? tag_input[21] : dirty_1_182; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3262 = waySel & _GEN_12323 ? tag_input[21] : dirty_1_183; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3263 = waySel & _GEN_12325 ? tag_input[21] : dirty_1_184; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3264 = waySel & _GEN_12327 ? tag_input[21] : dirty_1_185; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3265 = waySel & _GEN_12329 ? tag_input[21] : dirty_1_186; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3266 = waySel & _GEN_12331 ? tag_input[21] : dirty_1_187; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3267 = waySel & _GEN_12333 ? tag_input[21] : dirty_1_188; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3268 = waySel & _GEN_12335 ? tag_input[21] : dirty_1_189; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3269 = waySel & _GEN_12337 ? tag_input[21] : dirty_1_190; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3270 = waySel & _GEN_12339 ? tag_input[21] : dirty_1_191; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3271 = waySel & _GEN_12341 ? tag_input[21] : dirty_1_192; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3272 = waySel & _GEN_12343 ? tag_input[21] : dirty_1_193; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3273 = waySel & _GEN_12345 ? tag_input[21] : dirty_1_194; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3274 = waySel & _GEN_12347 ? tag_input[21] : dirty_1_195; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3275 = waySel & _GEN_12349 ? tag_input[21] : dirty_1_196; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3276 = waySel & _GEN_12351 ? tag_input[21] : dirty_1_197; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3277 = waySel & _GEN_12353 ? tag_input[21] : dirty_1_198; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3278 = waySel & _GEN_12355 ? tag_input[21] : dirty_1_199; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3279 = waySel & _GEN_12357 ? tag_input[21] : dirty_1_200; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3280 = waySel & _GEN_12359 ? tag_input[21] : dirty_1_201; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3281 = waySel & _GEN_12361 ? tag_input[21] : dirty_1_202; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3282 = waySel & _GEN_12363 ? tag_input[21] : dirty_1_203; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3283 = waySel & _GEN_12365 ? tag_input[21] : dirty_1_204; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3284 = waySel & _GEN_12367 ? tag_input[21] : dirty_1_205; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3285 = waySel & _GEN_12369 ? tag_input[21] : dirty_1_206; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3286 = waySel & _GEN_12371 ? tag_input[21] : dirty_1_207; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3287 = waySel & _GEN_12373 ? tag_input[21] : dirty_1_208; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3288 = waySel & _GEN_12375 ? tag_input[21] : dirty_1_209; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3289 = waySel & _GEN_12377 ? tag_input[21] : dirty_1_210; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3290 = waySel & _GEN_12379 ? tag_input[21] : dirty_1_211; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3291 = waySel & _GEN_12381 ? tag_input[21] : dirty_1_212; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3292 = waySel & _GEN_12383 ? tag_input[21] : dirty_1_213; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3293 = waySel & _GEN_12385 ? tag_input[21] : dirty_1_214; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3294 = waySel & _GEN_12387 ? tag_input[21] : dirty_1_215; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3295 = waySel & _GEN_12389 ? tag_input[21] : dirty_1_216; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3296 = waySel & _GEN_12391 ? tag_input[21] : dirty_1_217; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3297 = waySel & _GEN_12393 ? tag_input[21] : dirty_1_218; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3298 = waySel & _GEN_12395 ? tag_input[21] : dirty_1_219; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3299 = waySel & _GEN_12397 ? tag_input[21] : dirty_1_220; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3300 = waySel & _GEN_12399 ? tag_input[21] : dirty_1_221; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3301 = waySel & _GEN_12401 ? tag_input[21] : dirty_1_222; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3302 = waySel & _GEN_12403 ? tag_input[21] : dirty_1_223; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3303 = waySel & _GEN_12405 ? tag_input[21] : dirty_1_224; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3304 = waySel & _GEN_12407 ? tag_input[21] : dirty_1_225; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3305 = waySel & _GEN_12409 ? tag_input[21] : dirty_1_226; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3306 = waySel & _GEN_12411 ? tag_input[21] : dirty_1_227; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3307 = waySel & _GEN_12413 ? tag_input[21] : dirty_1_228; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3308 = waySel & _GEN_12415 ? tag_input[21] : dirty_1_229; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3309 = waySel & _GEN_12417 ? tag_input[21] : dirty_1_230; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3310 = waySel & _GEN_12419 ? tag_input[21] : dirty_1_231; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3311 = waySel & _GEN_12421 ? tag_input[21] : dirty_1_232; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3312 = waySel & _GEN_12423 ? tag_input[21] : dirty_1_233; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3313 = waySel & _GEN_12425 ? tag_input[21] : dirty_1_234; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3314 = waySel & _GEN_12427 ? tag_input[21] : dirty_1_235; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3315 = waySel & _GEN_12429 ? tag_input[21] : dirty_1_236; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3316 = waySel & _GEN_12431 ? tag_input[21] : dirty_1_237; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3317 = waySel & _GEN_12433 ? tag_input[21] : dirty_1_238; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3318 = waySel & _GEN_12435 ? tag_input[21] : dirty_1_239; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3319 = waySel & _GEN_12437 ? tag_input[21] : dirty_1_240; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3320 = waySel & _GEN_12439 ? tag_input[21] : dirty_1_241; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3321 = waySel & _GEN_12441 ? tag_input[21] : dirty_1_242; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3322 = waySel & _GEN_12443 ? tag_input[21] : dirty_1_243; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3323 = waySel & _GEN_12445 ? tag_input[21] : dirty_1_244; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3324 = waySel & _GEN_12447 ? tag_input[21] : dirty_1_245; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3325 = waySel & _GEN_12449 ? tag_input[21] : dirty_1_246; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3326 = waySel & _GEN_12451 ? tag_input[21] : dirty_1_247; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3327 = waySel & _GEN_12453 ? tag_input[21] : dirty_1_248; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3328 = waySel & _GEN_12455 ? tag_input[21] : dirty_1_249; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3329 = waySel & _GEN_12457 ? tag_input[21] : dirty_1_250; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3330 = waySel & _GEN_12459 ? tag_input[21] : dirty_1_251; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3331 = waySel & _GEN_12461 ? tag_input[21] : dirty_1_252; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3332 = waySel & _GEN_12463 ? tag_input[21] : dirty_1_253; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3333 = waySel & _GEN_12465 ? tag_input[21] : dirty_1_254; // @[dcache.scala 113:28 414:{66,66}]
  wire  _GEN_3334 = waySel & _GEN_12467 ? tag_input[21] : dirty_1_255; // @[dcache.scala 113:28 414:{66,66}]
  wire [20:0] _GEN_3335 = storeTag ? _GEN_2819 : 21'h0; // @[dcache.scala 143:25 411:31]
  wire [20:0] _GEN_3336 = storeTag ? _GEN_2820 : 21'h0; // @[dcache.scala 143:25 411:31]
  wire  _GEN_3337 = storeTag & _GEN_13518; // @[dcache.scala 144:25 411:31]
  wire  _GEN_3338 = storeTag & waySel; // @[dcache.scala 144:25 411:31]
  wire  _GEN_3339 = storeTag ? _GEN_2823 : dirty_0_0; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3340 = storeTag ? _GEN_2824 : dirty_0_1; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3341 = storeTag ? _GEN_2825 : dirty_0_2; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3342 = storeTag ? _GEN_2826 : dirty_0_3; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3343 = storeTag ? _GEN_2827 : dirty_0_4; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3344 = storeTag ? _GEN_2828 : dirty_0_5; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3345 = storeTag ? _GEN_2829 : dirty_0_6; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3346 = storeTag ? _GEN_2830 : dirty_0_7; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3347 = storeTag ? _GEN_2831 : dirty_0_8; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3348 = storeTag ? _GEN_2832 : dirty_0_9; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3349 = storeTag ? _GEN_2833 : dirty_0_10; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3350 = storeTag ? _GEN_2834 : dirty_0_11; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3351 = storeTag ? _GEN_2835 : dirty_0_12; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3352 = storeTag ? _GEN_2836 : dirty_0_13; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3353 = storeTag ? _GEN_2837 : dirty_0_14; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3354 = storeTag ? _GEN_2838 : dirty_0_15; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3355 = storeTag ? _GEN_2839 : dirty_0_16; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3356 = storeTag ? _GEN_2840 : dirty_0_17; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3357 = storeTag ? _GEN_2841 : dirty_0_18; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3358 = storeTag ? _GEN_2842 : dirty_0_19; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3359 = storeTag ? _GEN_2843 : dirty_0_20; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3360 = storeTag ? _GEN_2844 : dirty_0_21; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3361 = storeTag ? _GEN_2845 : dirty_0_22; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3362 = storeTag ? _GEN_2846 : dirty_0_23; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3363 = storeTag ? _GEN_2847 : dirty_0_24; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3364 = storeTag ? _GEN_2848 : dirty_0_25; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3365 = storeTag ? _GEN_2849 : dirty_0_26; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3366 = storeTag ? _GEN_2850 : dirty_0_27; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3367 = storeTag ? _GEN_2851 : dirty_0_28; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3368 = storeTag ? _GEN_2852 : dirty_0_29; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3369 = storeTag ? _GEN_2853 : dirty_0_30; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3370 = storeTag ? _GEN_2854 : dirty_0_31; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3371 = storeTag ? _GEN_2855 : dirty_0_32; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3372 = storeTag ? _GEN_2856 : dirty_0_33; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3373 = storeTag ? _GEN_2857 : dirty_0_34; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3374 = storeTag ? _GEN_2858 : dirty_0_35; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3375 = storeTag ? _GEN_2859 : dirty_0_36; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3376 = storeTag ? _GEN_2860 : dirty_0_37; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3377 = storeTag ? _GEN_2861 : dirty_0_38; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3378 = storeTag ? _GEN_2862 : dirty_0_39; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3379 = storeTag ? _GEN_2863 : dirty_0_40; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3380 = storeTag ? _GEN_2864 : dirty_0_41; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3381 = storeTag ? _GEN_2865 : dirty_0_42; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3382 = storeTag ? _GEN_2866 : dirty_0_43; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3383 = storeTag ? _GEN_2867 : dirty_0_44; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3384 = storeTag ? _GEN_2868 : dirty_0_45; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3385 = storeTag ? _GEN_2869 : dirty_0_46; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3386 = storeTag ? _GEN_2870 : dirty_0_47; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3387 = storeTag ? _GEN_2871 : dirty_0_48; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3388 = storeTag ? _GEN_2872 : dirty_0_49; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3389 = storeTag ? _GEN_2873 : dirty_0_50; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3390 = storeTag ? _GEN_2874 : dirty_0_51; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3391 = storeTag ? _GEN_2875 : dirty_0_52; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3392 = storeTag ? _GEN_2876 : dirty_0_53; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3393 = storeTag ? _GEN_2877 : dirty_0_54; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3394 = storeTag ? _GEN_2878 : dirty_0_55; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3395 = storeTag ? _GEN_2879 : dirty_0_56; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3396 = storeTag ? _GEN_2880 : dirty_0_57; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3397 = storeTag ? _GEN_2881 : dirty_0_58; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3398 = storeTag ? _GEN_2882 : dirty_0_59; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3399 = storeTag ? _GEN_2883 : dirty_0_60; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3400 = storeTag ? _GEN_2884 : dirty_0_61; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3401 = storeTag ? _GEN_2885 : dirty_0_62; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3402 = storeTag ? _GEN_2886 : dirty_0_63; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3403 = storeTag ? _GEN_2887 : dirty_0_64; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3404 = storeTag ? _GEN_2888 : dirty_0_65; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3405 = storeTag ? _GEN_2889 : dirty_0_66; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3406 = storeTag ? _GEN_2890 : dirty_0_67; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3407 = storeTag ? _GEN_2891 : dirty_0_68; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3408 = storeTag ? _GEN_2892 : dirty_0_69; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3409 = storeTag ? _GEN_2893 : dirty_0_70; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3410 = storeTag ? _GEN_2894 : dirty_0_71; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3411 = storeTag ? _GEN_2895 : dirty_0_72; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3412 = storeTag ? _GEN_2896 : dirty_0_73; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3413 = storeTag ? _GEN_2897 : dirty_0_74; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3414 = storeTag ? _GEN_2898 : dirty_0_75; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3415 = storeTag ? _GEN_2899 : dirty_0_76; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3416 = storeTag ? _GEN_2900 : dirty_0_77; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3417 = storeTag ? _GEN_2901 : dirty_0_78; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3418 = storeTag ? _GEN_2902 : dirty_0_79; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3419 = storeTag ? _GEN_2903 : dirty_0_80; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3420 = storeTag ? _GEN_2904 : dirty_0_81; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3421 = storeTag ? _GEN_2905 : dirty_0_82; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3422 = storeTag ? _GEN_2906 : dirty_0_83; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3423 = storeTag ? _GEN_2907 : dirty_0_84; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3424 = storeTag ? _GEN_2908 : dirty_0_85; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3425 = storeTag ? _GEN_2909 : dirty_0_86; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3426 = storeTag ? _GEN_2910 : dirty_0_87; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3427 = storeTag ? _GEN_2911 : dirty_0_88; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3428 = storeTag ? _GEN_2912 : dirty_0_89; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3429 = storeTag ? _GEN_2913 : dirty_0_90; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3430 = storeTag ? _GEN_2914 : dirty_0_91; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3431 = storeTag ? _GEN_2915 : dirty_0_92; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3432 = storeTag ? _GEN_2916 : dirty_0_93; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3433 = storeTag ? _GEN_2917 : dirty_0_94; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3434 = storeTag ? _GEN_2918 : dirty_0_95; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3435 = storeTag ? _GEN_2919 : dirty_0_96; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3436 = storeTag ? _GEN_2920 : dirty_0_97; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3437 = storeTag ? _GEN_2921 : dirty_0_98; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3438 = storeTag ? _GEN_2922 : dirty_0_99; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3439 = storeTag ? _GEN_2923 : dirty_0_100; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3440 = storeTag ? _GEN_2924 : dirty_0_101; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3441 = storeTag ? _GEN_2925 : dirty_0_102; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3442 = storeTag ? _GEN_2926 : dirty_0_103; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3443 = storeTag ? _GEN_2927 : dirty_0_104; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3444 = storeTag ? _GEN_2928 : dirty_0_105; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3445 = storeTag ? _GEN_2929 : dirty_0_106; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3446 = storeTag ? _GEN_2930 : dirty_0_107; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3447 = storeTag ? _GEN_2931 : dirty_0_108; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3448 = storeTag ? _GEN_2932 : dirty_0_109; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3449 = storeTag ? _GEN_2933 : dirty_0_110; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3450 = storeTag ? _GEN_2934 : dirty_0_111; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3451 = storeTag ? _GEN_2935 : dirty_0_112; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3452 = storeTag ? _GEN_2936 : dirty_0_113; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3453 = storeTag ? _GEN_2937 : dirty_0_114; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3454 = storeTag ? _GEN_2938 : dirty_0_115; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3455 = storeTag ? _GEN_2939 : dirty_0_116; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3456 = storeTag ? _GEN_2940 : dirty_0_117; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3457 = storeTag ? _GEN_2941 : dirty_0_118; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3458 = storeTag ? _GEN_2942 : dirty_0_119; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3459 = storeTag ? _GEN_2943 : dirty_0_120; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3460 = storeTag ? _GEN_2944 : dirty_0_121; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3461 = storeTag ? _GEN_2945 : dirty_0_122; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3462 = storeTag ? _GEN_2946 : dirty_0_123; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3463 = storeTag ? _GEN_2947 : dirty_0_124; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3464 = storeTag ? _GEN_2948 : dirty_0_125; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3465 = storeTag ? _GEN_2949 : dirty_0_126; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3466 = storeTag ? _GEN_2950 : dirty_0_127; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3467 = storeTag ? _GEN_2951 : dirty_0_128; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3468 = storeTag ? _GEN_2952 : dirty_0_129; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3469 = storeTag ? _GEN_2953 : dirty_0_130; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3470 = storeTag ? _GEN_2954 : dirty_0_131; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3471 = storeTag ? _GEN_2955 : dirty_0_132; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3472 = storeTag ? _GEN_2956 : dirty_0_133; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3473 = storeTag ? _GEN_2957 : dirty_0_134; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3474 = storeTag ? _GEN_2958 : dirty_0_135; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3475 = storeTag ? _GEN_2959 : dirty_0_136; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3476 = storeTag ? _GEN_2960 : dirty_0_137; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3477 = storeTag ? _GEN_2961 : dirty_0_138; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3478 = storeTag ? _GEN_2962 : dirty_0_139; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3479 = storeTag ? _GEN_2963 : dirty_0_140; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3480 = storeTag ? _GEN_2964 : dirty_0_141; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3481 = storeTag ? _GEN_2965 : dirty_0_142; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3482 = storeTag ? _GEN_2966 : dirty_0_143; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3483 = storeTag ? _GEN_2967 : dirty_0_144; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3484 = storeTag ? _GEN_2968 : dirty_0_145; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3485 = storeTag ? _GEN_2969 : dirty_0_146; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3486 = storeTag ? _GEN_2970 : dirty_0_147; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3487 = storeTag ? _GEN_2971 : dirty_0_148; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3488 = storeTag ? _GEN_2972 : dirty_0_149; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3489 = storeTag ? _GEN_2973 : dirty_0_150; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3490 = storeTag ? _GEN_2974 : dirty_0_151; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3491 = storeTag ? _GEN_2975 : dirty_0_152; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3492 = storeTag ? _GEN_2976 : dirty_0_153; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3493 = storeTag ? _GEN_2977 : dirty_0_154; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3494 = storeTag ? _GEN_2978 : dirty_0_155; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3495 = storeTag ? _GEN_2979 : dirty_0_156; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3496 = storeTag ? _GEN_2980 : dirty_0_157; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3497 = storeTag ? _GEN_2981 : dirty_0_158; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3498 = storeTag ? _GEN_2982 : dirty_0_159; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3499 = storeTag ? _GEN_2983 : dirty_0_160; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3500 = storeTag ? _GEN_2984 : dirty_0_161; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3501 = storeTag ? _GEN_2985 : dirty_0_162; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3502 = storeTag ? _GEN_2986 : dirty_0_163; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3503 = storeTag ? _GEN_2987 : dirty_0_164; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3504 = storeTag ? _GEN_2988 : dirty_0_165; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3505 = storeTag ? _GEN_2989 : dirty_0_166; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3506 = storeTag ? _GEN_2990 : dirty_0_167; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3507 = storeTag ? _GEN_2991 : dirty_0_168; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3508 = storeTag ? _GEN_2992 : dirty_0_169; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3509 = storeTag ? _GEN_2993 : dirty_0_170; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3510 = storeTag ? _GEN_2994 : dirty_0_171; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3511 = storeTag ? _GEN_2995 : dirty_0_172; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3512 = storeTag ? _GEN_2996 : dirty_0_173; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3513 = storeTag ? _GEN_2997 : dirty_0_174; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3514 = storeTag ? _GEN_2998 : dirty_0_175; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3515 = storeTag ? _GEN_2999 : dirty_0_176; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3516 = storeTag ? _GEN_3000 : dirty_0_177; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3517 = storeTag ? _GEN_3001 : dirty_0_178; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3518 = storeTag ? _GEN_3002 : dirty_0_179; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3519 = storeTag ? _GEN_3003 : dirty_0_180; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3520 = storeTag ? _GEN_3004 : dirty_0_181; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3521 = storeTag ? _GEN_3005 : dirty_0_182; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3522 = storeTag ? _GEN_3006 : dirty_0_183; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3523 = storeTag ? _GEN_3007 : dirty_0_184; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3524 = storeTag ? _GEN_3008 : dirty_0_185; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3525 = storeTag ? _GEN_3009 : dirty_0_186; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3526 = storeTag ? _GEN_3010 : dirty_0_187; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3527 = storeTag ? _GEN_3011 : dirty_0_188; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3528 = storeTag ? _GEN_3012 : dirty_0_189; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3529 = storeTag ? _GEN_3013 : dirty_0_190; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3530 = storeTag ? _GEN_3014 : dirty_0_191; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3531 = storeTag ? _GEN_3015 : dirty_0_192; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3532 = storeTag ? _GEN_3016 : dirty_0_193; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3533 = storeTag ? _GEN_3017 : dirty_0_194; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3534 = storeTag ? _GEN_3018 : dirty_0_195; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3535 = storeTag ? _GEN_3019 : dirty_0_196; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3536 = storeTag ? _GEN_3020 : dirty_0_197; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3537 = storeTag ? _GEN_3021 : dirty_0_198; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3538 = storeTag ? _GEN_3022 : dirty_0_199; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3539 = storeTag ? _GEN_3023 : dirty_0_200; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3540 = storeTag ? _GEN_3024 : dirty_0_201; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3541 = storeTag ? _GEN_3025 : dirty_0_202; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3542 = storeTag ? _GEN_3026 : dirty_0_203; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3543 = storeTag ? _GEN_3027 : dirty_0_204; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3544 = storeTag ? _GEN_3028 : dirty_0_205; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3545 = storeTag ? _GEN_3029 : dirty_0_206; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3546 = storeTag ? _GEN_3030 : dirty_0_207; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3547 = storeTag ? _GEN_3031 : dirty_0_208; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3548 = storeTag ? _GEN_3032 : dirty_0_209; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3549 = storeTag ? _GEN_3033 : dirty_0_210; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3550 = storeTag ? _GEN_3034 : dirty_0_211; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3551 = storeTag ? _GEN_3035 : dirty_0_212; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3552 = storeTag ? _GEN_3036 : dirty_0_213; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3553 = storeTag ? _GEN_3037 : dirty_0_214; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3554 = storeTag ? _GEN_3038 : dirty_0_215; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3555 = storeTag ? _GEN_3039 : dirty_0_216; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3556 = storeTag ? _GEN_3040 : dirty_0_217; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3557 = storeTag ? _GEN_3041 : dirty_0_218; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3558 = storeTag ? _GEN_3042 : dirty_0_219; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3559 = storeTag ? _GEN_3043 : dirty_0_220; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3560 = storeTag ? _GEN_3044 : dirty_0_221; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3561 = storeTag ? _GEN_3045 : dirty_0_222; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3562 = storeTag ? _GEN_3046 : dirty_0_223; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3563 = storeTag ? _GEN_3047 : dirty_0_224; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3564 = storeTag ? _GEN_3048 : dirty_0_225; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3565 = storeTag ? _GEN_3049 : dirty_0_226; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3566 = storeTag ? _GEN_3050 : dirty_0_227; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3567 = storeTag ? _GEN_3051 : dirty_0_228; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3568 = storeTag ? _GEN_3052 : dirty_0_229; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3569 = storeTag ? _GEN_3053 : dirty_0_230; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3570 = storeTag ? _GEN_3054 : dirty_0_231; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3571 = storeTag ? _GEN_3055 : dirty_0_232; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3572 = storeTag ? _GEN_3056 : dirty_0_233; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3573 = storeTag ? _GEN_3057 : dirty_0_234; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3574 = storeTag ? _GEN_3058 : dirty_0_235; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3575 = storeTag ? _GEN_3059 : dirty_0_236; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3576 = storeTag ? _GEN_3060 : dirty_0_237; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3577 = storeTag ? _GEN_3061 : dirty_0_238; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3578 = storeTag ? _GEN_3062 : dirty_0_239; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3579 = storeTag ? _GEN_3063 : dirty_0_240; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3580 = storeTag ? _GEN_3064 : dirty_0_241; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3581 = storeTag ? _GEN_3065 : dirty_0_242; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3582 = storeTag ? _GEN_3066 : dirty_0_243; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3583 = storeTag ? _GEN_3067 : dirty_0_244; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3584 = storeTag ? _GEN_3068 : dirty_0_245; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3585 = storeTag ? _GEN_3069 : dirty_0_246; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3586 = storeTag ? _GEN_3070 : dirty_0_247; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3587 = storeTag ? _GEN_3071 : dirty_0_248; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3588 = storeTag ? _GEN_3072 : dirty_0_249; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3589 = storeTag ? _GEN_3073 : dirty_0_250; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3590 = storeTag ? _GEN_3074 : dirty_0_251; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3591 = storeTag ? _GEN_3075 : dirty_0_252; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3592 = storeTag ? _GEN_3076 : dirty_0_253; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3593 = storeTag ? _GEN_3077 : dirty_0_254; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3594 = storeTag ? _GEN_3078 : dirty_0_255; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3595 = storeTag ? _GEN_3079 : dirty_1_0; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3596 = storeTag ? _GEN_3080 : dirty_1_1; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3597 = storeTag ? _GEN_3081 : dirty_1_2; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3598 = storeTag ? _GEN_3082 : dirty_1_3; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3599 = storeTag ? _GEN_3083 : dirty_1_4; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3600 = storeTag ? _GEN_3084 : dirty_1_5; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3601 = storeTag ? _GEN_3085 : dirty_1_6; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3602 = storeTag ? _GEN_3086 : dirty_1_7; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3603 = storeTag ? _GEN_3087 : dirty_1_8; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3604 = storeTag ? _GEN_3088 : dirty_1_9; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3605 = storeTag ? _GEN_3089 : dirty_1_10; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3606 = storeTag ? _GEN_3090 : dirty_1_11; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3607 = storeTag ? _GEN_3091 : dirty_1_12; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3608 = storeTag ? _GEN_3092 : dirty_1_13; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3609 = storeTag ? _GEN_3093 : dirty_1_14; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3610 = storeTag ? _GEN_3094 : dirty_1_15; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3611 = storeTag ? _GEN_3095 : dirty_1_16; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3612 = storeTag ? _GEN_3096 : dirty_1_17; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3613 = storeTag ? _GEN_3097 : dirty_1_18; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3614 = storeTag ? _GEN_3098 : dirty_1_19; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3615 = storeTag ? _GEN_3099 : dirty_1_20; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3616 = storeTag ? _GEN_3100 : dirty_1_21; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3617 = storeTag ? _GEN_3101 : dirty_1_22; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3618 = storeTag ? _GEN_3102 : dirty_1_23; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3619 = storeTag ? _GEN_3103 : dirty_1_24; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3620 = storeTag ? _GEN_3104 : dirty_1_25; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3621 = storeTag ? _GEN_3105 : dirty_1_26; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3622 = storeTag ? _GEN_3106 : dirty_1_27; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3623 = storeTag ? _GEN_3107 : dirty_1_28; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3624 = storeTag ? _GEN_3108 : dirty_1_29; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3625 = storeTag ? _GEN_3109 : dirty_1_30; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3626 = storeTag ? _GEN_3110 : dirty_1_31; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3627 = storeTag ? _GEN_3111 : dirty_1_32; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3628 = storeTag ? _GEN_3112 : dirty_1_33; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3629 = storeTag ? _GEN_3113 : dirty_1_34; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3630 = storeTag ? _GEN_3114 : dirty_1_35; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3631 = storeTag ? _GEN_3115 : dirty_1_36; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3632 = storeTag ? _GEN_3116 : dirty_1_37; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3633 = storeTag ? _GEN_3117 : dirty_1_38; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3634 = storeTag ? _GEN_3118 : dirty_1_39; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3635 = storeTag ? _GEN_3119 : dirty_1_40; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3636 = storeTag ? _GEN_3120 : dirty_1_41; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3637 = storeTag ? _GEN_3121 : dirty_1_42; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3638 = storeTag ? _GEN_3122 : dirty_1_43; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3639 = storeTag ? _GEN_3123 : dirty_1_44; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3640 = storeTag ? _GEN_3124 : dirty_1_45; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3641 = storeTag ? _GEN_3125 : dirty_1_46; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3642 = storeTag ? _GEN_3126 : dirty_1_47; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3643 = storeTag ? _GEN_3127 : dirty_1_48; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3644 = storeTag ? _GEN_3128 : dirty_1_49; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3645 = storeTag ? _GEN_3129 : dirty_1_50; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3646 = storeTag ? _GEN_3130 : dirty_1_51; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3647 = storeTag ? _GEN_3131 : dirty_1_52; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3648 = storeTag ? _GEN_3132 : dirty_1_53; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3649 = storeTag ? _GEN_3133 : dirty_1_54; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3650 = storeTag ? _GEN_3134 : dirty_1_55; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3651 = storeTag ? _GEN_3135 : dirty_1_56; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3652 = storeTag ? _GEN_3136 : dirty_1_57; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3653 = storeTag ? _GEN_3137 : dirty_1_58; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3654 = storeTag ? _GEN_3138 : dirty_1_59; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3655 = storeTag ? _GEN_3139 : dirty_1_60; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3656 = storeTag ? _GEN_3140 : dirty_1_61; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3657 = storeTag ? _GEN_3141 : dirty_1_62; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3658 = storeTag ? _GEN_3142 : dirty_1_63; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3659 = storeTag ? _GEN_3143 : dirty_1_64; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3660 = storeTag ? _GEN_3144 : dirty_1_65; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3661 = storeTag ? _GEN_3145 : dirty_1_66; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3662 = storeTag ? _GEN_3146 : dirty_1_67; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3663 = storeTag ? _GEN_3147 : dirty_1_68; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3664 = storeTag ? _GEN_3148 : dirty_1_69; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3665 = storeTag ? _GEN_3149 : dirty_1_70; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3666 = storeTag ? _GEN_3150 : dirty_1_71; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3667 = storeTag ? _GEN_3151 : dirty_1_72; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3668 = storeTag ? _GEN_3152 : dirty_1_73; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3669 = storeTag ? _GEN_3153 : dirty_1_74; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3670 = storeTag ? _GEN_3154 : dirty_1_75; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3671 = storeTag ? _GEN_3155 : dirty_1_76; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3672 = storeTag ? _GEN_3156 : dirty_1_77; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3673 = storeTag ? _GEN_3157 : dirty_1_78; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3674 = storeTag ? _GEN_3158 : dirty_1_79; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3675 = storeTag ? _GEN_3159 : dirty_1_80; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3676 = storeTag ? _GEN_3160 : dirty_1_81; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3677 = storeTag ? _GEN_3161 : dirty_1_82; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3678 = storeTag ? _GEN_3162 : dirty_1_83; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3679 = storeTag ? _GEN_3163 : dirty_1_84; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3680 = storeTag ? _GEN_3164 : dirty_1_85; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3681 = storeTag ? _GEN_3165 : dirty_1_86; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3682 = storeTag ? _GEN_3166 : dirty_1_87; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3683 = storeTag ? _GEN_3167 : dirty_1_88; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3684 = storeTag ? _GEN_3168 : dirty_1_89; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3685 = storeTag ? _GEN_3169 : dirty_1_90; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3686 = storeTag ? _GEN_3170 : dirty_1_91; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3687 = storeTag ? _GEN_3171 : dirty_1_92; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3688 = storeTag ? _GEN_3172 : dirty_1_93; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3689 = storeTag ? _GEN_3173 : dirty_1_94; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3690 = storeTag ? _GEN_3174 : dirty_1_95; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3691 = storeTag ? _GEN_3175 : dirty_1_96; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3692 = storeTag ? _GEN_3176 : dirty_1_97; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3693 = storeTag ? _GEN_3177 : dirty_1_98; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3694 = storeTag ? _GEN_3178 : dirty_1_99; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3695 = storeTag ? _GEN_3179 : dirty_1_100; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3696 = storeTag ? _GEN_3180 : dirty_1_101; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3697 = storeTag ? _GEN_3181 : dirty_1_102; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3698 = storeTag ? _GEN_3182 : dirty_1_103; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3699 = storeTag ? _GEN_3183 : dirty_1_104; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3700 = storeTag ? _GEN_3184 : dirty_1_105; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3701 = storeTag ? _GEN_3185 : dirty_1_106; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3702 = storeTag ? _GEN_3186 : dirty_1_107; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3703 = storeTag ? _GEN_3187 : dirty_1_108; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3704 = storeTag ? _GEN_3188 : dirty_1_109; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3705 = storeTag ? _GEN_3189 : dirty_1_110; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3706 = storeTag ? _GEN_3190 : dirty_1_111; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3707 = storeTag ? _GEN_3191 : dirty_1_112; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3708 = storeTag ? _GEN_3192 : dirty_1_113; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3709 = storeTag ? _GEN_3193 : dirty_1_114; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3710 = storeTag ? _GEN_3194 : dirty_1_115; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3711 = storeTag ? _GEN_3195 : dirty_1_116; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3712 = storeTag ? _GEN_3196 : dirty_1_117; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3713 = storeTag ? _GEN_3197 : dirty_1_118; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3714 = storeTag ? _GEN_3198 : dirty_1_119; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3715 = storeTag ? _GEN_3199 : dirty_1_120; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3716 = storeTag ? _GEN_3200 : dirty_1_121; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3717 = storeTag ? _GEN_3201 : dirty_1_122; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3718 = storeTag ? _GEN_3202 : dirty_1_123; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3719 = storeTag ? _GEN_3203 : dirty_1_124; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3720 = storeTag ? _GEN_3204 : dirty_1_125; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3721 = storeTag ? _GEN_3205 : dirty_1_126; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3722 = storeTag ? _GEN_3206 : dirty_1_127; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3723 = storeTag ? _GEN_3207 : dirty_1_128; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3724 = storeTag ? _GEN_3208 : dirty_1_129; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3725 = storeTag ? _GEN_3209 : dirty_1_130; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3726 = storeTag ? _GEN_3210 : dirty_1_131; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3727 = storeTag ? _GEN_3211 : dirty_1_132; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3728 = storeTag ? _GEN_3212 : dirty_1_133; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3729 = storeTag ? _GEN_3213 : dirty_1_134; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3730 = storeTag ? _GEN_3214 : dirty_1_135; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3731 = storeTag ? _GEN_3215 : dirty_1_136; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3732 = storeTag ? _GEN_3216 : dirty_1_137; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3733 = storeTag ? _GEN_3217 : dirty_1_138; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3734 = storeTag ? _GEN_3218 : dirty_1_139; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3735 = storeTag ? _GEN_3219 : dirty_1_140; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3736 = storeTag ? _GEN_3220 : dirty_1_141; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3737 = storeTag ? _GEN_3221 : dirty_1_142; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3738 = storeTag ? _GEN_3222 : dirty_1_143; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3739 = storeTag ? _GEN_3223 : dirty_1_144; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3740 = storeTag ? _GEN_3224 : dirty_1_145; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3741 = storeTag ? _GEN_3225 : dirty_1_146; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3742 = storeTag ? _GEN_3226 : dirty_1_147; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3743 = storeTag ? _GEN_3227 : dirty_1_148; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3744 = storeTag ? _GEN_3228 : dirty_1_149; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3745 = storeTag ? _GEN_3229 : dirty_1_150; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3746 = storeTag ? _GEN_3230 : dirty_1_151; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3747 = storeTag ? _GEN_3231 : dirty_1_152; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3748 = storeTag ? _GEN_3232 : dirty_1_153; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3749 = storeTag ? _GEN_3233 : dirty_1_154; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3750 = storeTag ? _GEN_3234 : dirty_1_155; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3751 = storeTag ? _GEN_3235 : dirty_1_156; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3752 = storeTag ? _GEN_3236 : dirty_1_157; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3753 = storeTag ? _GEN_3237 : dirty_1_158; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3754 = storeTag ? _GEN_3238 : dirty_1_159; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3755 = storeTag ? _GEN_3239 : dirty_1_160; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3756 = storeTag ? _GEN_3240 : dirty_1_161; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3757 = storeTag ? _GEN_3241 : dirty_1_162; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3758 = storeTag ? _GEN_3242 : dirty_1_163; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3759 = storeTag ? _GEN_3243 : dirty_1_164; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3760 = storeTag ? _GEN_3244 : dirty_1_165; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3761 = storeTag ? _GEN_3245 : dirty_1_166; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3762 = storeTag ? _GEN_3246 : dirty_1_167; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3763 = storeTag ? _GEN_3247 : dirty_1_168; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3764 = storeTag ? _GEN_3248 : dirty_1_169; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3765 = storeTag ? _GEN_3249 : dirty_1_170; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3766 = storeTag ? _GEN_3250 : dirty_1_171; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3767 = storeTag ? _GEN_3251 : dirty_1_172; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3768 = storeTag ? _GEN_3252 : dirty_1_173; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3769 = storeTag ? _GEN_3253 : dirty_1_174; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3770 = storeTag ? _GEN_3254 : dirty_1_175; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3771 = storeTag ? _GEN_3255 : dirty_1_176; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3772 = storeTag ? _GEN_3256 : dirty_1_177; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3773 = storeTag ? _GEN_3257 : dirty_1_178; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3774 = storeTag ? _GEN_3258 : dirty_1_179; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3775 = storeTag ? _GEN_3259 : dirty_1_180; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3776 = storeTag ? _GEN_3260 : dirty_1_181; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3777 = storeTag ? _GEN_3261 : dirty_1_182; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3778 = storeTag ? _GEN_3262 : dirty_1_183; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3779 = storeTag ? _GEN_3263 : dirty_1_184; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3780 = storeTag ? _GEN_3264 : dirty_1_185; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3781 = storeTag ? _GEN_3265 : dirty_1_186; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3782 = storeTag ? _GEN_3266 : dirty_1_187; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3783 = storeTag ? _GEN_3267 : dirty_1_188; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3784 = storeTag ? _GEN_3268 : dirty_1_189; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3785 = storeTag ? _GEN_3269 : dirty_1_190; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3786 = storeTag ? _GEN_3270 : dirty_1_191; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3787 = storeTag ? _GEN_3271 : dirty_1_192; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3788 = storeTag ? _GEN_3272 : dirty_1_193; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3789 = storeTag ? _GEN_3273 : dirty_1_194; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3790 = storeTag ? _GEN_3274 : dirty_1_195; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3791 = storeTag ? _GEN_3275 : dirty_1_196; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3792 = storeTag ? _GEN_3276 : dirty_1_197; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3793 = storeTag ? _GEN_3277 : dirty_1_198; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3794 = storeTag ? _GEN_3278 : dirty_1_199; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3795 = storeTag ? _GEN_3279 : dirty_1_200; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3796 = storeTag ? _GEN_3280 : dirty_1_201; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3797 = storeTag ? _GEN_3281 : dirty_1_202; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3798 = storeTag ? _GEN_3282 : dirty_1_203; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3799 = storeTag ? _GEN_3283 : dirty_1_204; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3800 = storeTag ? _GEN_3284 : dirty_1_205; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3801 = storeTag ? _GEN_3285 : dirty_1_206; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3802 = storeTag ? _GEN_3286 : dirty_1_207; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3803 = storeTag ? _GEN_3287 : dirty_1_208; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3804 = storeTag ? _GEN_3288 : dirty_1_209; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3805 = storeTag ? _GEN_3289 : dirty_1_210; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3806 = storeTag ? _GEN_3290 : dirty_1_211; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3807 = storeTag ? _GEN_3291 : dirty_1_212; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3808 = storeTag ? _GEN_3292 : dirty_1_213; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3809 = storeTag ? _GEN_3293 : dirty_1_214; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3810 = storeTag ? _GEN_3294 : dirty_1_215; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3811 = storeTag ? _GEN_3295 : dirty_1_216; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3812 = storeTag ? _GEN_3296 : dirty_1_217; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3813 = storeTag ? _GEN_3297 : dirty_1_218; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3814 = storeTag ? _GEN_3298 : dirty_1_219; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3815 = storeTag ? _GEN_3299 : dirty_1_220; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3816 = storeTag ? _GEN_3300 : dirty_1_221; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3817 = storeTag ? _GEN_3301 : dirty_1_222; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3818 = storeTag ? _GEN_3302 : dirty_1_223; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3819 = storeTag ? _GEN_3303 : dirty_1_224; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3820 = storeTag ? _GEN_3304 : dirty_1_225; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3821 = storeTag ? _GEN_3305 : dirty_1_226; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3822 = storeTag ? _GEN_3306 : dirty_1_227; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3823 = storeTag ? _GEN_3307 : dirty_1_228; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3824 = storeTag ? _GEN_3308 : dirty_1_229; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3825 = storeTag ? _GEN_3309 : dirty_1_230; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3826 = storeTag ? _GEN_3310 : dirty_1_231; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3827 = storeTag ? _GEN_3311 : dirty_1_232; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3828 = storeTag ? _GEN_3312 : dirty_1_233; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3829 = storeTag ? _GEN_3313 : dirty_1_234; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3830 = storeTag ? _GEN_3314 : dirty_1_235; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3831 = storeTag ? _GEN_3315 : dirty_1_236; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3832 = storeTag ? _GEN_3316 : dirty_1_237; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3833 = storeTag ? _GEN_3317 : dirty_1_238; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3834 = storeTag ? _GEN_3318 : dirty_1_239; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3835 = storeTag ? _GEN_3319 : dirty_1_240; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3836 = storeTag ? _GEN_3320 : dirty_1_241; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3837 = storeTag ? _GEN_3321 : dirty_1_242; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3838 = storeTag ? _GEN_3322 : dirty_1_243; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3839 = storeTag ? _GEN_3323 : dirty_1_244; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3840 = storeTag ? _GEN_3324 : dirty_1_245; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3841 = storeTag ? _GEN_3325 : dirty_1_246; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3842 = storeTag ? _GEN_3326 : dirty_1_247; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3843 = storeTag ? _GEN_3327 : dirty_1_248; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3844 = storeTag ? _GEN_3328 : dirty_1_249; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3845 = storeTag ? _GEN_3329 : dirty_1_250; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3846 = storeTag ? _GEN_3330 : dirty_1_251; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3847 = storeTag ? _GEN_3331 : dirty_1_252; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3848 = storeTag ? _GEN_3332 : dirty_1_253; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3849 = storeTag ? _GEN_3333 : dirty_1_254; // @[dcache.scala 113:28 411:31]
  wire  _GEN_3850 = storeTag ? _GEN_3334 : dirty_1_255; // @[dcache.scala 113:28 411:31]
  wire [20:0] _GEN_3851 = ~waySel ? 21'h0 : _GEN_3335; // @[dcache.scala 418:{66,66}]
  wire [20:0] _GEN_3852 = waySel ? 21'h0 : _GEN_3336; // @[dcache.scala 418:{66,66}]
  wire  _GEN_3853 = _GEN_13518 | _GEN_3337; // @[dcache.scala 419:{66,66}]
  wire  _GEN_3854 = waySel | _GEN_3338; // @[dcache.scala 419:{66,66}]
  wire  _GEN_3855 = _GEN_13518 & _GEN_12468 ? 1'h0 : _GEN_3339; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3856 = _GEN_13518 & _GEN_11959 ? 1'h0 : _GEN_3340; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3857 = _GEN_13518 & _GEN_11961 ? 1'h0 : _GEN_3341; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3858 = _GEN_13518 & _GEN_11963 ? 1'h0 : _GEN_3342; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3859 = _GEN_13518 & _GEN_11965 ? 1'h0 : _GEN_3343; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3860 = _GEN_13518 & _GEN_11967 ? 1'h0 : _GEN_3344; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3861 = _GEN_13518 & _GEN_11969 ? 1'h0 : _GEN_3345; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3862 = _GEN_13518 & _GEN_11971 ? 1'h0 : _GEN_3346; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3863 = _GEN_13518 & _GEN_11973 ? 1'h0 : _GEN_3347; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3864 = _GEN_13518 & _GEN_11975 ? 1'h0 : _GEN_3348; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3865 = _GEN_13518 & _GEN_11977 ? 1'h0 : _GEN_3349; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3866 = _GEN_13518 & _GEN_11979 ? 1'h0 : _GEN_3350; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3867 = _GEN_13518 & _GEN_11981 ? 1'h0 : _GEN_3351; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3868 = _GEN_13518 & _GEN_11983 ? 1'h0 : _GEN_3352; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3869 = _GEN_13518 & _GEN_11985 ? 1'h0 : _GEN_3353; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3870 = _GEN_13518 & _GEN_11987 ? 1'h0 : _GEN_3354; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3871 = _GEN_13518 & _GEN_11989 ? 1'h0 : _GEN_3355; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3872 = _GEN_13518 & _GEN_11991 ? 1'h0 : _GEN_3356; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3873 = _GEN_13518 & _GEN_11993 ? 1'h0 : _GEN_3357; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3874 = _GEN_13518 & _GEN_11995 ? 1'h0 : _GEN_3358; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3875 = _GEN_13518 & _GEN_11997 ? 1'h0 : _GEN_3359; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3876 = _GEN_13518 & _GEN_11999 ? 1'h0 : _GEN_3360; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3877 = _GEN_13518 & _GEN_12001 ? 1'h0 : _GEN_3361; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3878 = _GEN_13518 & _GEN_12003 ? 1'h0 : _GEN_3362; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3879 = _GEN_13518 & _GEN_12005 ? 1'h0 : _GEN_3363; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3880 = _GEN_13518 & _GEN_12007 ? 1'h0 : _GEN_3364; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3881 = _GEN_13518 & _GEN_12009 ? 1'h0 : _GEN_3365; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3882 = _GEN_13518 & _GEN_12011 ? 1'h0 : _GEN_3366; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3883 = _GEN_13518 & _GEN_12013 ? 1'h0 : _GEN_3367; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3884 = _GEN_13518 & _GEN_12015 ? 1'h0 : _GEN_3368; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3885 = _GEN_13518 & _GEN_12017 ? 1'h0 : _GEN_3369; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3886 = _GEN_13518 & _GEN_12019 ? 1'h0 : _GEN_3370; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3887 = _GEN_13518 & _GEN_12021 ? 1'h0 : _GEN_3371; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3888 = _GEN_13518 & _GEN_12023 ? 1'h0 : _GEN_3372; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3889 = _GEN_13518 & _GEN_12025 ? 1'h0 : _GEN_3373; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3890 = _GEN_13518 & _GEN_12027 ? 1'h0 : _GEN_3374; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3891 = _GEN_13518 & _GEN_12029 ? 1'h0 : _GEN_3375; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3892 = _GEN_13518 & _GEN_12031 ? 1'h0 : _GEN_3376; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3893 = _GEN_13518 & _GEN_12033 ? 1'h0 : _GEN_3377; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3894 = _GEN_13518 & _GEN_12035 ? 1'h0 : _GEN_3378; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3895 = _GEN_13518 & _GEN_12037 ? 1'h0 : _GEN_3379; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3896 = _GEN_13518 & _GEN_12039 ? 1'h0 : _GEN_3380; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3897 = _GEN_13518 & _GEN_12041 ? 1'h0 : _GEN_3381; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3898 = _GEN_13518 & _GEN_12043 ? 1'h0 : _GEN_3382; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3899 = _GEN_13518 & _GEN_12045 ? 1'h0 : _GEN_3383; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3900 = _GEN_13518 & _GEN_12047 ? 1'h0 : _GEN_3384; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3901 = _GEN_13518 & _GEN_12049 ? 1'h0 : _GEN_3385; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3902 = _GEN_13518 & _GEN_12051 ? 1'h0 : _GEN_3386; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3903 = _GEN_13518 & _GEN_12053 ? 1'h0 : _GEN_3387; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3904 = _GEN_13518 & _GEN_12055 ? 1'h0 : _GEN_3388; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3905 = _GEN_13518 & _GEN_12057 ? 1'h0 : _GEN_3389; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3906 = _GEN_13518 & _GEN_12059 ? 1'h0 : _GEN_3390; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3907 = _GEN_13518 & _GEN_12061 ? 1'h0 : _GEN_3391; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3908 = _GEN_13518 & _GEN_12063 ? 1'h0 : _GEN_3392; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3909 = _GEN_13518 & _GEN_12065 ? 1'h0 : _GEN_3393; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3910 = _GEN_13518 & _GEN_12067 ? 1'h0 : _GEN_3394; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3911 = _GEN_13518 & _GEN_12069 ? 1'h0 : _GEN_3395; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3912 = _GEN_13518 & _GEN_12071 ? 1'h0 : _GEN_3396; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3913 = _GEN_13518 & _GEN_12073 ? 1'h0 : _GEN_3397; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3914 = _GEN_13518 & _GEN_12075 ? 1'h0 : _GEN_3398; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3915 = _GEN_13518 & _GEN_12077 ? 1'h0 : _GEN_3399; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3916 = _GEN_13518 & _GEN_12079 ? 1'h0 : _GEN_3400; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3917 = _GEN_13518 & _GEN_12081 ? 1'h0 : _GEN_3401; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3918 = _GEN_13518 & _GEN_12083 ? 1'h0 : _GEN_3402; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3919 = _GEN_13518 & _GEN_12085 ? 1'h0 : _GEN_3403; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3920 = _GEN_13518 & _GEN_12087 ? 1'h0 : _GEN_3404; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3921 = _GEN_13518 & _GEN_12089 ? 1'h0 : _GEN_3405; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3922 = _GEN_13518 & _GEN_12091 ? 1'h0 : _GEN_3406; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3923 = _GEN_13518 & _GEN_12093 ? 1'h0 : _GEN_3407; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3924 = _GEN_13518 & _GEN_12095 ? 1'h0 : _GEN_3408; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3925 = _GEN_13518 & _GEN_12097 ? 1'h0 : _GEN_3409; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3926 = _GEN_13518 & _GEN_12099 ? 1'h0 : _GEN_3410; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3927 = _GEN_13518 & _GEN_12101 ? 1'h0 : _GEN_3411; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3928 = _GEN_13518 & _GEN_12103 ? 1'h0 : _GEN_3412; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3929 = _GEN_13518 & _GEN_12105 ? 1'h0 : _GEN_3413; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3930 = _GEN_13518 & _GEN_12107 ? 1'h0 : _GEN_3414; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3931 = _GEN_13518 & _GEN_12109 ? 1'h0 : _GEN_3415; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3932 = _GEN_13518 & _GEN_12111 ? 1'h0 : _GEN_3416; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3933 = _GEN_13518 & _GEN_12113 ? 1'h0 : _GEN_3417; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3934 = _GEN_13518 & _GEN_12115 ? 1'h0 : _GEN_3418; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3935 = _GEN_13518 & _GEN_12117 ? 1'h0 : _GEN_3419; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3936 = _GEN_13518 & _GEN_12119 ? 1'h0 : _GEN_3420; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3937 = _GEN_13518 & _GEN_12121 ? 1'h0 : _GEN_3421; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3938 = _GEN_13518 & _GEN_12123 ? 1'h0 : _GEN_3422; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3939 = _GEN_13518 & _GEN_12125 ? 1'h0 : _GEN_3423; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3940 = _GEN_13518 & _GEN_12127 ? 1'h0 : _GEN_3424; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3941 = _GEN_13518 & _GEN_12129 ? 1'h0 : _GEN_3425; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3942 = _GEN_13518 & _GEN_12131 ? 1'h0 : _GEN_3426; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3943 = _GEN_13518 & _GEN_12133 ? 1'h0 : _GEN_3427; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3944 = _GEN_13518 & _GEN_12135 ? 1'h0 : _GEN_3428; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3945 = _GEN_13518 & _GEN_12137 ? 1'h0 : _GEN_3429; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3946 = _GEN_13518 & _GEN_12139 ? 1'h0 : _GEN_3430; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3947 = _GEN_13518 & _GEN_12141 ? 1'h0 : _GEN_3431; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3948 = _GEN_13518 & _GEN_12143 ? 1'h0 : _GEN_3432; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3949 = _GEN_13518 & _GEN_12145 ? 1'h0 : _GEN_3433; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3950 = _GEN_13518 & _GEN_12147 ? 1'h0 : _GEN_3434; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3951 = _GEN_13518 & _GEN_12149 ? 1'h0 : _GEN_3435; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3952 = _GEN_13518 & _GEN_12151 ? 1'h0 : _GEN_3436; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3953 = _GEN_13518 & _GEN_12153 ? 1'h0 : _GEN_3437; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3954 = _GEN_13518 & _GEN_12155 ? 1'h0 : _GEN_3438; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3955 = _GEN_13518 & _GEN_12157 ? 1'h0 : _GEN_3439; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3956 = _GEN_13518 & _GEN_12159 ? 1'h0 : _GEN_3440; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3957 = _GEN_13518 & _GEN_12161 ? 1'h0 : _GEN_3441; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3958 = _GEN_13518 & _GEN_12163 ? 1'h0 : _GEN_3442; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3959 = _GEN_13518 & _GEN_12165 ? 1'h0 : _GEN_3443; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3960 = _GEN_13518 & _GEN_12167 ? 1'h0 : _GEN_3444; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3961 = _GEN_13518 & _GEN_12169 ? 1'h0 : _GEN_3445; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3962 = _GEN_13518 & _GEN_12171 ? 1'h0 : _GEN_3446; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3963 = _GEN_13518 & _GEN_12173 ? 1'h0 : _GEN_3447; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3964 = _GEN_13518 & _GEN_12175 ? 1'h0 : _GEN_3448; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3965 = _GEN_13518 & _GEN_12177 ? 1'h0 : _GEN_3449; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3966 = _GEN_13518 & _GEN_12179 ? 1'h0 : _GEN_3450; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3967 = _GEN_13518 & _GEN_12181 ? 1'h0 : _GEN_3451; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3968 = _GEN_13518 & _GEN_12183 ? 1'h0 : _GEN_3452; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3969 = _GEN_13518 & _GEN_12185 ? 1'h0 : _GEN_3453; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3970 = _GEN_13518 & _GEN_12187 ? 1'h0 : _GEN_3454; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3971 = _GEN_13518 & _GEN_12189 ? 1'h0 : _GEN_3455; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3972 = _GEN_13518 & _GEN_12191 ? 1'h0 : _GEN_3456; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3973 = _GEN_13518 & _GEN_12193 ? 1'h0 : _GEN_3457; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3974 = _GEN_13518 & _GEN_12195 ? 1'h0 : _GEN_3458; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3975 = _GEN_13518 & _GEN_12197 ? 1'h0 : _GEN_3459; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3976 = _GEN_13518 & _GEN_12199 ? 1'h0 : _GEN_3460; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3977 = _GEN_13518 & _GEN_12201 ? 1'h0 : _GEN_3461; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3978 = _GEN_13518 & _GEN_12203 ? 1'h0 : _GEN_3462; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3979 = _GEN_13518 & _GEN_12205 ? 1'h0 : _GEN_3463; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3980 = _GEN_13518 & _GEN_12207 ? 1'h0 : _GEN_3464; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3981 = _GEN_13518 & _GEN_12209 ? 1'h0 : _GEN_3465; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3982 = _GEN_13518 & _GEN_12211 ? 1'h0 : _GEN_3466; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3983 = _GEN_13518 & _GEN_12213 ? 1'h0 : _GEN_3467; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3984 = _GEN_13518 & _GEN_12215 ? 1'h0 : _GEN_3468; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3985 = _GEN_13518 & _GEN_12217 ? 1'h0 : _GEN_3469; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3986 = _GEN_13518 & _GEN_12219 ? 1'h0 : _GEN_3470; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3987 = _GEN_13518 & _GEN_12221 ? 1'h0 : _GEN_3471; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3988 = _GEN_13518 & _GEN_12223 ? 1'h0 : _GEN_3472; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3989 = _GEN_13518 & _GEN_12225 ? 1'h0 : _GEN_3473; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3990 = _GEN_13518 & _GEN_12227 ? 1'h0 : _GEN_3474; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3991 = _GEN_13518 & _GEN_12229 ? 1'h0 : _GEN_3475; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3992 = _GEN_13518 & _GEN_12231 ? 1'h0 : _GEN_3476; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3993 = _GEN_13518 & _GEN_12233 ? 1'h0 : _GEN_3477; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3994 = _GEN_13518 & _GEN_12235 ? 1'h0 : _GEN_3478; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3995 = _GEN_13518 & _GEN_12237 ? 1'h0 : _GEN_3479; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3996 = _GEN_13518 & _GEN_12239 ? 1'h0 : _GEN_3480; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3997 = _GEN_13518 & _GEN_12241 ? 1'h0 : _GEN_3481; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3998 = _GEN_13518 & _GEN_12243 ? 1'h0 : _GEN_3482; // @[dcache.scala 420:{66,66}]
  wire  _GEN_3999 = _GEN_13518 & _GEN_12245 ? 1'h0 : _GEN_3483; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4000 = _GEN_13518 & _GEN_12247 ? 1'h0 : _GEN_3484; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4001 = _GEN_13518 & _GEN_12249 ? 1'h0 : _GEN_3485; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4002 = _GEN_13518 & _GEN_12251 ? 1'h0 : _GEN_3486; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4003 = _GEN_13518 & _GEN_12253 ? 1'h0 : _GEN_3487; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4004 = _GEN_13518 & _GEN_12255 ? 1'h0 : _GEN_3488; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4005 = _GEN_13518 & _GEN_12257 ? 1'h0 : _GEN_3489; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4006 = _GEN_13518 & _GEN_12259 ? 1'h0 : _GEN_3490; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4007 = _GEN_13518 & _GEN_12261 ? 1'h0 : _GEN_3491; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4008 = _GEN_13518 & _GEN_12263 ? 1'h0 : _GEN_3492; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4009 = _GEN_13518 & _GEN_12265 ? 1'h0 : _GEN_3493; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4010 = _GEN_13518 & _GEN_12267 ? 1'h0 : _GEN_3494; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4011 = _GEN_13518 & _GEN_12269 ? 1'h0 : _GEN_3495; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4012 = _GEN_13518 & _GEN_12271 ? 1'h0 : _GEN_3496; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4013 = _GEN_13518 & _GEN_12273 ? 1'h0 : _GEN_3497; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4014 = _GEN_13518 & _GEN_12275 ? 1'h0 : _GEN_3498; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4015 = _GEN_13518 & _GEN_12277 ? 1'h0 : _GEN_3499; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4016 = _GEN_13518 & _GEN_12279 ? 1'h0 : _GEN_3500; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4017 = _GEN_13518 & _GEN_12281 ? 1'h0 : _GEN_3501; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4018 = _GEN_13518 & _GEN_12283 ? 1'h0 : _GEN_3502; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4019 = _GEN_13518 & _GEN_12285 ? 1'h0 : _GEN_3503; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4020 = _GEN_13518 & _GEN_12287 ? 1'h0 : _GEN_3504; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4021 = _GEN_13518 & _GEN_12289 ? 1'h0 : _GEN_3505; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4022 = _GEN_13518 & _GEN_12291 ? 1'h0 : _GEN_3506; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4023 = _GEN_13518 & _GEN_12293 ? 1'h0 : _GEN_3507; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4024 = _GEN_13518 & _GEN_12295 ? 1'h0 : _GEN_3508; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4025 = _GEN_13518 & _GEN_12297 ? 1'h0 : _GEN_3509; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4026 = _GEN_13518 & _GEN_12299 ? 1'h0 : _GEN_3510; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4027 = _GEN_13518 & _GEN_12301 ? 1'h0 : _GEN_3511; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4028 = _GEN_13518 & _GEN_12303 ? 1'h0 : _GEN_3512; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4029 = _GEN_13518 & _GEN_12305 ? 1'h0 : _GEN_3513; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4030 = _GEN_13518 & _GEN_12307 ? 1'h0 : _GEN_3514; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4031 = _GEN_13518 & _GEN_12309 ? 1'h0 : _GEN_3515; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4032 = _GEN_13518 & _GEN_12311 ? 1'h0 : _GEN_3516; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4033 = _GEN_13518 & _GEN_12313 ? 1'h0 : _GEN_3517; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4034 = _GEN_13518 & _GEN_12315 ? 1'h0 : _GEN_3518; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4035 = _GEN_13518 & _GEN_12317 ? 1'h0 : _GEN_3519; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4036 = _GEN_13518 & _GEN_12319 ? 1'h0 : _GEN_3520; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4037 = _GEN_13518 & _GEN_12321 ? 1'h0 : _GEN_3521; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4038 = _GEN_13518 & _GEN_12323 ? 1'h0 : _GEN_3522; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4039 = _GEN_13518 & _GEN_12325 ? 1'h0 : _GEN_3523; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4040 = _GEN_13518 & _GEN_12327 ? 1'h0 : _GEN_3524; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4041 = _GEN_13518 & _GEN_12329 ? 1'h0 : _GEN_3525; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4042 = _GEN_13518 & _GEN_12331 ? 1'h0 : _GEN_3526; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4043 = _GEN_13518 & _GEN_12333 ? 1'h0 : _GEN_3527; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4044 = _GEN_13518 & _GEN_12335 ? 1'h0 : _GEN_3528; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4045 = _GEN_13518 & _GEN_12337 ? 1'h0 : _GEN_3529; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4046 = _GEN_13518 & _GEN_12339 ? 1'h0 : _GEN_3530; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4047 = _GEN_13518 & _GEN_12341 ? 1'h0 : _GEN_3531; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4048 = _GEN_13518 & _GEN_12343 ? 1'h0 : _GEN_3532; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4049 = _GEN_13518 & _GEN_12345 ? 1'h0 : _GEN_3533; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4050 = _GEN_13518 & _GEN_12347 ? 1'h0 : _GEN_3534; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4051 = _GEN_13518 & _GEN_12349 ? 1'h0 : _GEN_3535; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4052 = _GEN_13518 & _GEN_12351 ? 1'h0 : _GEN_3536; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4053 = _GEN_13518 & _GEN_12353 ? 1'h0 : _GEN_3537; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4054 = _GEN_13518 & _GEN_12355 ? 1'h0 : _GEN_3538; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4055 = _GEN_13518 & _GEN_12357 ? 1'h0 : _GEN_3539; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4056 = _GEN_13518 & _GEN_12359 ? 1'h0 : _GEN_3540; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4057 = _GEN_13518 & _GEN_12361 ? 1'h0 : _GEN_3541; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4058 = _GEN_13518 & _GEN_12363 ? 1'h0 : _GEN_3542; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4059 = _GEN_13518 & _GEN_12365 ? 1'h0 : _GEN_3543; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4060 = _GEN_13518 & _GEN_12367 ? 1'h0 : _GEN_3544; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4061 = _GEN_13518 & _GEN_12369 ? 1'h0 : _GEN_3545; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4062 = _GEN_13518 & _GEN_12371 ? 1'h0 : _GEN_3546; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4063 = _GEN_13518 & _GEN_12373 ? 1'h0 : _GEN_3547; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4064 = _GEN_13518 & _GEN_12375 ? 1'h0 : _GEN_3548; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4065 = _GEN_13518 & _GEN_12377 ? 1'h0 : _GEN_3549; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4066 = _GEN_13518 & _GEN_12379 ? 1'h0 : _GEN_3550; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4067 = _GEN_13518 & _GEN_12381 ? 1'h0 : _GEN_3551; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4068 = _GEN_13518 & _GEN_12383 ? 1'h0 : _GEN_3552; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4069 = _GEN_13518 & _GEN_12385 ? 1'h0 : _GEN_3553; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4070 = _GEN_13518 & _GEN_12387 ? 1'h0 : _GEN_3554; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4071 = _GEN_13518 & _GEN_12389 ? 1'h0 : _GEN_3555; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4072 = _GEN_13518 & _GEN_12391 ? 1'h0 : _GEN_3556; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4073 = _GEN_13518 & _GEN_12393 ? 1'h0 : _GEN_3557; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4074 = _GEN_13518 & _GEN_12395 ? 1'h0 : _GEN_3558; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4075 = _GEN_13518 & _GEN_12397 ? 1'h0 : _GEN_3559; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4076 = _GEN_13518 & _GEN_12399 ? 1'h0 : _GEN_3560; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4077 = _GEN_13518 & _GEN_12401 ? 1'h0 : _GEN_3561; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4078 = _GEN_13518 & _GEN_12403 ? 1'h0 : _GEN_3562; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4079 = _GEN_13518 & _GEN_12405 ? 1'h0 : _GEN_3563; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4080 = _GEN_13518 & _GEN_12407 ? 1'h0 : _GEN_3564; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4081 = _GEN_13518 & _GEN_12409 ? 1'h0 : _GEN_3565; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4082 = _GEN_13518 & _GEN_12411 ? 1'h0 : _GEN_3566; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4083 = _GEN_13518 & _GEN_12413 ? 1'h0 : _GEN_3567; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4084 = _GEN_13518 & _GEN_12415 ? 1'h0 : _GEN_3568; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4085 = _GEN_13518 & _GEN_12417 ? 1'h0 : _GEN_3569; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4086 = _GEN_13518 & _GEN_12419 ? 1'h0 : _GEN_3570; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4087 = _GEN_13518 & _GEN_12421 ? 1'h0 : _GEN_3571; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4088 = _GEN_13518 & _GEN_12423 ? 1'h0 : _GEN_3572; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4089 = _GEN_13518 & _GEN_12425 ? 1'h0 : _GEN_3573; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4090 = _GEN_13518 & _GEN_12427 ? 1'h0 : _GEN_3574; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4091 = _GEN_13518 & _GEN_12429 ? 1'h0 : _GEN_3575; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4092 = _GEN_13518 & _GEN_12431 ? 1'h0 : _GEN_3576; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4093 = _GEN_13518 & _GEN_12433 ? 1'h0 : _GEN_3577; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4094 = _GEN_13518 & _GEN_12435 ? 1'h0 : _GEN_3578; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4095 = _GEN_13518 & _GEN_12437 ? 1'h0 : _GEN_3579; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4096 = _GEN_13518 & _GEN_12439 ? 1'h0 : _GEN_3580; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4097 = _GEN_13518 & _GEN_12441 ? 1'h0 : _GEN_3581; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4098 = _GEN_13518 & _GEN_12443 ? 1'h0 : _GEN_3582; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4099 = _GEN_13518 & _GEN_12445 ? 1'h0 : _GEN_3583; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4100 = _GEN_13518 & _GEN_12447 ? 1'h0 : _GEN_3584; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4101 = _GEN_13518 & _GEN_12449 ? 1'h0 : _GEN_3585; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4102 = _GEN_13518 & _GEN_12451 ? 1'h0 : _GEN_3586; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4103 = _GEN_13518 & _GEN_12453 ? 1'h0 : _GEN_3587; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4104 = _GEN_13518 & _GEN_12455 ? 1'h0 : _GEN_3588; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4105 = _GEN_13518 & _GEN_12457 ? 1'h0 : _GEN_3589; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4106 = _GEN_13518 & _GEN_12459 ? 1'h0 : _GEN_3590; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4107 = _GEN_13518 & _GEN_12461 ? 1'h0 : _GEN_3591; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4108 = _GEN_13518 & _GEN_12463 ? 1'h0 : _GEN_3592; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4109 = _GEN_13518 & _GEN_12465 ? 1'h0 : _GEN_3593; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4110 = _GEN_13518 & _GEN_12467 ? 1'h0 : _GEN_3594; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4111 = waySel & _GEN_12468 ? 1'h0 : _GEN_3595; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4112 = waySel & _GEN_11959 ? 1'h0 : _GEN_3596; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4113 = waySel & _GEN_11961 ? 1'h0 : _GEN_3597; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4114 = waySel & _GEN_11963 ? 1'h0 : _GEN_3598; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4115 = waySel & _GEN_11965 ? 1'h0 : _GEN_3599; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4116 = waySel & _GEN_11967 ? 1'h0 : _GEN_3600; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4117 = waySel & _GEN_11969 ? 1'h0 : _GEN_3601; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4118 = waySel & _GEN_11971 ? 1'h0 : _GEN_3602; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4119 = waySel & _GEN_11973 ? 1'h0 : _GEN_3603; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4120 = waySel & _GEN_11975 ? 1'h0 : _GEN_3604; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4121 = waySel & _GEN_11977 ? 1'h0 : _GEN_3605; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4122 = waySel & _GEN_11979 ? 1'h0 : _GEN_3606; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4123 = waySel & _GEN_11981 ? 1'h0 : _GEN_3607; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4124 = waySel & _GEN_11983 ? 1'h0 : _GEN_3608; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4125 = waySel & _GEN_11985 ? 1'h0 : _GEN_3609; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4126 = waySel & _GEN_11987 ? 1'h0 : _GEN_3610; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4127 = waySel & _GEN_11989 ? 1'h0 : _GEN_3611; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4128 = waySel & _GEN_11991 ? 1'h0 : _GEN_3612; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4129 = waySel & _GEN_11993 ? 1'h0 : _GEN_3613; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4130 = waySel & _GEN_11995 ? 1'h0 : _GEN_3614; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4131 = waySel & _GEN_11997 ? 1'h0 : _GEN_3615; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4132 = waySel & _GEN_11999 ? 1'h0 : _GEN_3616; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4133 = waySel & _GEN_12001 ? 1'h0 : _GEN_3617; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4134 = waySel & _GEN_12003 ? 1'h0 : _GEN_3618; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4135 = waySel & _GEN_12005 ? 1'h0 : _GEN_3619; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4136 = waySel & _GEN_12007 ? 1'h0 : _GEN_3620; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4137 = waySel & _GEN_12009 ? 1'h0 : _GEN_3621; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4138 = waySel & _GEN_12011 ? 1'h0 : _GEN_3622; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4139 = waySel & _GEN_12013 ? 1'h0 : _GEN_3623; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4140 = waySel & _GEN_12015 ? 1'h0 : _GEN_3624; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4141 = waySel & _GEN_12017 ? 1'h0 : _GEN_3625; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4142 = waySel & _GEN_12019 ? 1'h0 : _GEN_3626; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4143 = waySel & _GEN_12021 ? 1'h0 : _GEN_3627; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4144 = waySel & _GEN_12023 ? 1'h0 : _GEN_3628; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4145 = waySel & _GEN_12025 ? 1'h0 : _GEN_3629; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4146 = waySel & _GEN_12027 ? 1'h0 : _GEN_3630; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4147 = waySel & _GEN_12029 ? 1'h0 : _GEN_3631; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4148 = waySel & _GEN_12031 ? 1'h0 : _GEN_3632; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4149 = waySel & _GEN_12033 ? 1'h0 : _GEN_3633; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4150 = waySel & _GEN_12035 ? 1'h0 : _GEN_3634; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4151 = waySel & _GEN_12037 ? 1'h0 : _GEN_3635; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4152 = waySel & _GEN_12039 ? 1'h0 : _GEN_3636; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4153 = waySel & _GEN_12041 ? 1'h0 : _GEN_3637; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4154 = waySel & _GEN_12043 ? 1'h0 : _GEN_3638; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4155 = waySel & _GEN_12045 ? 1'h0 : _GEN_3639; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4156 = waySel & _GEN_12047 ? 1'h0 : _GEN_3640; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4157 = waySel & _GEN_12049 ? 1'h0 : _GEN_3641; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4158 = waySel & _GEN_12051 ? 1'h0 : _GEN_3642; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4159 = waySel & _GEN_12053 ? 1'h0 : _GEN_3643; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4160 = waySel & _GEN_12055 ? 1'h0 : _GEN_3644; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4161 = waySel & _GEN_12057 ? 1'h0 : _GEN_3645; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4162 = waySel & _GEN_12059 ? 1'h0 : _GEN_3646; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4163 = waySel & _GEN_12061 ? 1'h0 : _GEN_3647; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4164 = waySel & _GEN_12063 ? 1'h0 : _GEN_3648; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4165 = waySel & _GEN_12065 ? 1'h0 : _GEN_3649; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4166 = waySel & _GEN_12067 ? 1'h0 : _GEN_3650; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4167 = waySel & _GEN_12069 ? 1'h0 : _GEN_3651; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4168 = waySel & _GEN_12071 ? 1'h0 : _GEN_3652; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4169 = waySel & _GEN_12073 ? 1'h0 : _GEN_3653; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4170 = waySel & _GEN_12075 ? 1'h0 : _GEN_3654; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4171 = waySel & _GEN_12077 ? 1'h0 : _GEN_3655; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4172 = waySel & _GEN_12079 ? 1'h0 : _GEN_3656; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4173 = waySel & _GEN_12081 ? 1'h0 : _GEN_3657; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4174 = waySel & _GEN_12083 ? 1'h0 : _GEN_3658; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4175 = waySel & _GEN_12085 ? 1'h0 : _GEN_3659; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4176 = waySel & _GEN_12087 ? 1'h0 : _GEN_3660; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4177 = waySel & _GEN_12089 ? 1'h0 : _GEN_3661; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4178 = waySel & _GEN_12091 ? 1'h0 : _GEN_3662; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4179 = waySel & _GEN_12093 ? 1'h0 : _GEN_3663; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4180 = waySel & _GEN_12095 ? 1'h0 : _GEN_3664; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4181 = waySel & _GEN_12097 ? 1'h0 : _GEN_3665; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4182 = waySel & _GEN_12099 ? 1'h0 : _GEN_3666; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4183 = waySel & _GEN_12101 ? 1'h0 : _GEN_3667; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4184 = waySel & _GEN_12103 ? 1'h0 : _GEN_3668; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4185 = waySel & _GEN_12105 ? 1'h0 : _GEN_3669; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4186 = waySel & _GEN_12107 ? 1'h0 : _GEN_3670; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4187 = waySel & _GEN_12109 ? 1'h0 : _GEN_3671; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4188 = waySel & _GEN_12111 ? 1'h0 : _GEN_3672; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4189 = waySel & _GEN_12113 ? 1'h0 : _GEN_3673; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4190 = waySel & _GEN_12115 ? 1'h0 : _GEN_3674; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4191 = waySel & _GEN_12117 ? 1'h0 : _GEN_3675; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4192 = waySel & _GEN_12119 ? 1'h0 : _GEN_3676; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4193 = waySel & _GEN_12121 ? 1'h0 : _GEN_3677; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4194 = waySel & _GEN_12123 ? 1'h0 : _GEN_3678; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4195 = waySel & _GEN_12125 ? 1'h0 : _GEN_3679; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4196 = waySel & _GEN_12127 ? 1'h0 : _GEN_3680; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4197 = waySel & _GEN_12129 ? 1'h0 : _GEN_3681; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4198 = waySel & _GEN_12131 ? 1'h0 : _GEN_3682; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4199 = waySel & _GEN_12133 ? 1'h0 : _GEN_3683; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4200 = waySel & _GEN_12135 ? 1'h0 : _GEN_3684; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4201 = waySel & _GEN_12137 ? 1'h0 : _GEN_3685; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4202 = waySel & _GEN_12139 ? 1'h0 : _GEN_3686; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4203 = waySel & _GEN_12141 ? 1'h0 : _GEN_3687; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4204 = waySel & _GEN_12143 ? 1'h0 : _GEN_3688; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4205 = waySel & _GEN_12145 ? 1'h0 : _GEN_3689; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4206 = waySel & _GEN_12147 ? 1'h0 : _GEN_3690; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4207 = waySel & _GEN_12149 ? 1'h0 : _GEN_3691; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4208 = waySel & _GEN_12151 ? 1'h0 : _GEN_3692; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4209 = waySel & _GEN_12153 ? 1'h0 : _GEN_3693; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4210 = waySel & _GEN_12155 ? 1'h0 : _GEN_3694; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4211 = waySel & _GEN_12157 ? 1'h0 : _GEN_3695; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4212 = waySel & _GEN_12159 ? 1'h0 : _GEN_3696; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4213 = waySel & _GEN_12161 ? 1'h0 : _GEN_3697; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4214 = waySel & _GEN_12163 ? 1'h0 : _GEN_3698; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4215 = waySel & _GEN_12165 ? 1'h0 : _GEN_3699; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4216 = waySel & _GEN_12167 ? 1'h0 : _GEN_3700; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4217 = waySel & _GEN_12169 ? 1'h0 : _GEN_3701; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4218 = waySel & _GEN_12171 ? 1'h0 : _GEN_3702; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4219 = waySel & _GEN_12173 ? 1'h0 : _GEN_3703; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4220 = waySel & _GEN_12175 ? 1'h0 : _GEN_3704; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4221 = waySel & _GEN_12177 ? 1'h0 : _GEN_3705; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4222 = waySel & _GEN_12179 ? 1'h0 : _GEN_3706; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4223 = waySel & _GEN_12181 ? 1'h0 : _GEN_3707; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4224 = waySel & _GEN_12183 ? 1'h0 : _GEN_3708; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4225 = waySel & _GEN_12185 ? 1'h0 : _GEN_3709; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4226 = waySel & _GEN_12187 ? 1'h0 : _GEN_3710; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4227 = waySel & _GEN_12189 ? 1'h0 : _GEN_3711; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4228 = waySel & _GEN_12191 ? 1'h0 : _GEN_3712; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4229 = waySel & _GEN_12193 ? 1'h0 : _GEN_3713; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4230 = waySel & _GEN_12195 ? 1'h0 : _GEN_3714; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4231 = waySel & _GEN_12197 ? 1'h0 : _GEN_3715; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4232 = waySel & _GEN_12199 ? 1'h0 : _GEN_3716; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4233 = waySel & _GEN_12201 ? 1'h0 : _GEN_3717; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4234 = waySel & _GEN_12203 ? 1'h0 : _GEN_3718; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4235 = waySel & _GEN_12205 ? 1'h0 : _GEN_3719; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4236 = waySel & _GEN_12207 ? 1'h0 : _GEN_3720; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4237 = waySel & _GEN_12209 ? 1'h0 : _GEN_3721; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4238 = waySel & _GEN_12211 ? 1'h0 : _GEN_3722; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4239 = waySel & _GEN_12213 ? 1'h0 : _GEN_3723; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4240 = waySel & _GEN_12215 ? 1'h0 : _GEN_3724; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4241 = waySel & _GEN_12217 ? 1'h0 : _GEN_3725; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4242 = waySel & _GEN_12219 ? 1'h0 : _GEN_3726; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4243 = waySel & _GEN_12221 ? 1'h0 : _GEN_3727; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4244 = waySel & _GEN_12223 ? 1'h0 : _GEN_3728; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4245 = waySel & _GEN_12225 ? 1'h0 : _GEN_3729; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4246 = waySel & _GEN_12227 ? 1'h0 : _GEN_3730; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4247 = waySel & _GEN_12229 ? 1'h0 : _GEN_3731; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4248 = waySel & _GEN_12231 ? 1'h0 : _GEN_3732; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4249 = waySel & _GEN_12233 ? 1'h0 : _GEN_3733; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4250 = waySel & _GEN_12235 ? 1'h0 : _GEN_3734; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4251 = waySel & _GEN_12237 ? 1'h0 : _GEN_3735; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4252 = waySel & _GEN_12239 ? 1'h0 : _GEN_3736; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4253 = waySel & _GEN_12241 ? 1'h0 : _GEN_3737; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4254 = waySel & _GEN_12243 ? 1'h0 : _GEN_3738; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4255 = waySel & _GEN_12245 ? 1'h0 : _GEN_3739; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4256 = waySel & _GEN_12247 ? 1'h0 : _GEN_3740; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4257 = waySel & _GEN_12249 ? 1'h0 : _GEN_3741; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4258 = waySel & _GEN_12251 ? 1'h0 : _GEN_3742; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4259 = waySel & _GEN_12253 ? 1'h0 : _GEN_3743; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4260 = waySel & _GEN_12255 ? 1'h0 : _GEN_3744; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4261 = waySel & _GEN_12257 ? 1'h0 : _GEN_3745; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4262 = waySel & _GEN_12259 ? 1'h0 : _GEN_3746; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4263 = waySel & _GEN_12261 ? 1'h0 : _GEN_3747; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4264 = waySel & _GEN_12263 ? 1'h0 : _GEN_3748; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4265 = waySel & _GEN_12265 ? 1'h0 : _GEN_3749; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4266 = waySel & _GEN_12267 ? 1'h0 : _GEN_3750; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4267 = waySel & _GEN_12269 ? 1'h0 : _GEN_3751; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4268 = waySel & _GEN_12271 ? 1'h0 : _GEN_3752; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4269 = waySel & _GEN_12273 ? 1'h0 : _GEN_3753; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4270 = waySel & _GEN_12275 ? 1'h0 : _GEN_3754; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4271 = waySel & _GEN_12277 ? 1'h0 : _GEN_3755; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4272 = waySel & _GEN_12279 ? 1'h0 : _GEN_3756; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4273 = waySel & _GEN_12281 ? 1'h0 : _GEN_3757; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4274 = waySel & _GEN_12283 ? 1'h0 : _GEN_3758; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4275 = waySel & _GEN_12285 ? 1'h0 : _GEN_3759; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4276 = waySel & _GEN_12287 ? 1'h0 : _GEN_3760; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4277 = waySel & _GEN_12289 ? 1'h0 : _GEN_3761; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4278 = waySel & _GEN_12291 ? 1'h0 : _GEN_3762; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4279 = waySel & _GEN_12293 ? 1'h0 : _GEN_3763; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4280 = waySel & _GEN_12295 ? 1'h0 : _GEN_3764; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4281 = waySel & _GEN_12297 ? 1'h0 : _GEN_3765; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4282 = waySel & _GEN_12299 ? 1'h0 : _GEN_3766; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4283 = waySel & _GEN_12301 ? 1'h0 : _GEN_3767; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4284 = waySel & _GEN_12303 ? 1'h0 : _GEN_3768; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4285 = waySel & _GEN_12305 ? 1'h0 : _GEN_3769; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4286 = waySel & _GEN_12307 ? 1'h0 : _GEN_3770; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4287 = waySel & _GEN_12309 ? 1'h0 : _GEN_3771; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4288 = waySel & _GEN_12311 ? 1'h0 : _GEN_3772; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4289 = waySel & _GEN_12313 ? 1'h0 : _GEN_3773; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4290 = waySel & _GEN_12315 ? 1'h0 : _GEN_3774; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4291 = waySel & _GEN_12317 ? 1'h0 : _GEN_3775; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4292 = waySel & _GEN_12319 ? 1'h0 : _GEN_3776; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4293 = waySel & _GEN_12321 ? 1'h0 : _GEN_3777; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4294 = waySel & _GEN_12323 ? 1'h0 : _GEN_3778; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4295 = waySel & _GEN_12325 ? 1'h0 : _GEN_3779; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4296 = waySel & _GEN_12327 ? 1'h0 : _GEN_3780; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4297 = waySel & _GEN_12329 ? 1'h0 : _GEN_3781; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4298 = waySel & _GEN_12331 ? 1'h0 : _GEN_3782; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4299 = waySel & _GEN_12333 ? 1'h0 : _GEN_3783; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4300 = waySel & _GEN_12335 ? 1'h0 : _GEN_3784; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4301 = waySel & _GEN_12337 ? 1'h0 : _GEN_3785; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4302 = waySel & _GEN_12339 ? 1'h0 : _GEN_3786; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4303 = waySel & _GEN_12341 ? 1'h0 : _GEN_3787; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4304 = waySel & _GEN_12343 ? 1'h0 : _GEN_3788; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4305 = waySel & _GEN_12345 ? 1'h0 : _GEN_3789; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4306 = waySel & _GEN_12347 ? 1'h0 : _GEN_3790; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4307 = waySel & _GEN_12349 ? 1'h0 : _GEN_3791; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4308 = waySel & _GEN_12351 ? 1'h0 : _GEN_3792; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4309 = waySel & _GEN_12353 ? 1'h0 : _GEN_3793; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4310 = waySel & _GEN_12355 ? 1'h0 : _GEN_3794; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4311 = waySel & _GEN_12357 ? 1'h0 : _GEN_3795; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4312 = waySel & _GEN_12359 ? 1'h0 : _GEN_3796; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4313 = waySel & _GEN_12361 ? 1'h0 : _GEN_3797; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4314 = waySel & _GEN_12363 ? 1'h0 : _GEN_3798; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4315 = waySel & _GEN_12365 ? 1'h0 : _GEN_3799; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4316 = waySel & _GEN_12367 ? 1'h0 : _GEN_3800; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4317 = waySel & _GEN_12369 ? 1'h0 : _GEN_3801; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4318 = waySel & _GEN_12371 ? 1'h0 : _GEN_3802; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4319 = waySel & _GEN_12373 ? 1'h0 : _GEN_3803; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4320 = waySel & _GEN_12375 ? 1'h0 : _GEN_3804; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4321 = waySel & _GEN_12377 ? 1'h0 : _GEN_3805; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4322 = waySel & _GEN_12379 ? 1'h0 : _GEN_3806; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4323 = waySel & _GEN_12381 ? 1'h0 : _GEN_3807; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4324 = waySel & _GEN_12383 ? 1'h0 : _GEN_3808; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4325 = waySel & _GEN_12385 ? 1'h0 : _GEN_3809; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4326 = waySel & _GEN_12387 ? 1'h0 : _GEN_3810; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4327 = waySel & _GEN_12389 ? 1'h0 : _GEN_3811; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4328 = waySel & _GEN_12391 ? 1'h0 : _GEN_3812; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4329 = waySel & _GEN_12393 ? 1'h0 : _GEN_3813; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4330 = waySel & _GEN_12395 ? 1'h0 : _GEN_3814; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4331 = waySel & _GEN_12397 ? 1'h0 : _GEN_3815; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4332 = waySel & _GEN_12399 ? 1'h0 : _GEN_3816; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4333 = waySel & _GEN_12401 ? 1'h0 : _GEN_3817; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4334 = waySel & _GEN_12403 ? 1'h0 : _GEN_3818; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4335 = waySel & _GEN_12405 ? 1'h0 : _GEN_3819; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4336 = waySel & _GEN_12407 ? 1'h0 : _GEN_3820; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4337 = waySel & _GEN_12409 ? 1'h0 : _GEN_3821; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4338 = waySel & _GEN_12411 ? 1'h0 : _GEN_3822; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4339 = waySel & _GEN_12413 ? 1'h0 : _GEN_3823; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4340 = waySel & _GEN_12415 ? 1'h0 : _GEN_3824; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4341 = waySel & _GEN_12417 ? 1'h0 : _GEN_3825; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4342 = waySel & _GEN_12419 ? 1'h0 : _GEN_3826; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4343 = waySel & _GEN_12421 ? 1'h0 : _GEN_3827; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4344 = waySel & _GEN_12423 ? 1'h0 : _GEN_3828; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4345 = waySel & _GEN_12425 ? 1'h0 : _GEN_3829; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4346 = waySel & _GEN_12427 ? 1'h0 : _GEN_3830; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4347 = waySel & _GEN_12429 ? 1'h0 : _GEN_3831; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4348 = waySel & _GEN_12431 ? 1'h0 : _GEN_3832; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4349 = waySel & _GEN_12433 ? 1'h0 : _GEN_3833; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4350 = waySel & _GEN_12435 ? 1'h0 : _GEN_3834; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4351 = waySel & _GEN_12437 ? 1'h0 : _GEN_3835; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4352 = waySel & _GEN_12439 ? 1'h0 : _GEN_3836; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4353 = waySel & _GEN_12441 ? 1'h0 : _GEN_3837; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4354 = waySel & _GEN_12443 ? 1'h0 : _GEN_3838; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4355 = waySel & _GEN_12445 ? 1'h0 : _GEN_3839; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4356 = waySel & _GEN_12447 ? 1'h0 : _GEN_3840; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4357 = waySel & _GEN_12449 ? 1'h0 : _GEN_3841; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4358 = waySel & _GEN_12451 ? 1'h0 : _GEN_3842; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4359 = waySel & _GEN_12453 ? 1'h0 : _GEN_3843; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4360 = waySel & _GEN_12455 ? 1'h0 : _GEN_3844; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4361 = waySel & _GEN_12457 ? 1'h0 : _GEN_3845; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4362 = waySel & _GEN_12459 ? 1'h0 : _GEN_3846; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4363 = waySel & _GEN_12461 ? 1'h0 : _GEN_3847; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4364 = waySel & _GEN_12463 ? 1'h0 : _GEN_3848; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4365 = waySel & _GEN_12465 ? 1'h0 : _GEN_3849; // @[dcache.scala 420:{66,66}]
  wire  _GEN_4366 = waySel & _GEN_12467 ? 1'h0 : _GEN_3850; // @[dcache.scala 420:{66,66}]
  wire [20:0] _GEN_4367 = ~refillIDX_r ? 21'h0 : _GEN_3335; // @[dcache.scala 422:{61,61}]
  wire [20:0] _GEN_4368 = refillIDX_r ? 21'h0 : _GEN_3336; // @[dcache.scala 422:{61,61}]
  wire  _GEN_4369 = _GEN_11958 | _GEN_3337; // @[dcache.scala 423:{61,61}]
  wire  _GEN_4370 = refillIDX_r | _GEN_3338; // @[dcache.scala 423:{61,61}]
  wire  _GEN_4371 = _GEN_11958 & _GEN_12468 ? 1'h0 : _GEN_3339; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4372 = _GEN_11958 & _GEN_11959 ? 1'h0 : _GEN_3340; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4373 = _GEN_11958 & _GEN_11961 ? 1'h0 : _GEN_3341; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4374 = _GEN_11958 & _GEN_11963 ? 1'h0 : _GEN_3342; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4375 = _GEN_11958 & _GEN_11965 ? 1'h0 : _GEN_3343; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4376 = _GEN_11958 & _GEN_11967 ? 1'h0 : _GEN_3344; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4377 = _GEN_11958 & _GEN_11969 ? 1'h0 : _GEN_3345; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4378 = _GEN_11958 & _GEN_11971 ? 1'h0 : _GEN_3346; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4379 = _GEN_11958 & _GEN_11973 ? 1'h0 : _GEN_3347; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4380 = _GEN_11958 & _GEN_11975 ? 1'h0 : _GEN_3348; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4381 = _GEN_11958 & _GEN_11977 ? 1'h0 : _GEN_3349; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4382 = _GEN_11958 & _GEN_11979 ? 1'h0 : _GEN_3350; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4383 = _GEN_11958 & _GEN_11981 ? 1'h0 : _GEN_3351; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4384 = _GEN_11958 & _GEN_11983 ? 1'h0 : _GEN_3352; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4385 = _GEN_11958 & _GEN_11985 ? 1'h0 : _GEN_3353; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4386 = _GEN_11958 & _GEN_11987 ? 1'h0 : _GEN_3354; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4387 = _GEN_11958 & _GEN_11989 ? 1'h0 : _GEN_3355; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4388 = _GEN_11958 & _GEN_11991 ? 1'h0 : _GEN_3356; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4389 = _GEN_11958 & _GEN_11993 ? 1'h0 : _GEN_3357; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4390 = _GEN_11958 & _GEN_11995 ? 1'h0 : _GEN_3358; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4391 = _GEN_11958 & _GEN_11997 ? 1'h0 : _GEN_3359; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4392 = _GEN_11958 & _GEN_11999 ? 1'h0 : _GEN_3360; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4393 = _GEN_11958 & _GEN_12001 ? 1'h0 : _GEN_3361; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4394 = _GEN_11958 & _GEN_12003 ? 1'h0 : _GEN_3362; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4395 = _GEN_11958 & _GEN_12005 ? 1'h0 : _GEN_3363; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4396 = _GEN_11958 & _GEN_12007 ? 1'h0 : _GEN_3364; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4397 = _GEN_11958 & _GEN_12009 ? 1'h0 : _GEN_3365; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4398 = _GEN_11958 & _GEN_12011 ? 1'h0 : _GEN_3366; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4399 = _GEN_11958 & _GEN_12013 ? 1'h0 : _GEN_3367; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4400 = _GEN_11958 & _GEN_12015 ? 1'h0 : _GEN_3368; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4401 = _GEN_11958 & _GEN_12017 ? 1'h0 : _GEN_3369; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4402 = _GEN_11958 & _GEN_12019 ? 1'h0 : _GEN_3370; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4403 = _GEN_11958 & _GEN_12021 ? 1'h0 : _GEN_3371; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4404 = _GEN_11958 & _GEN_12023 ? 1'h0 : _GEN_3372; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4405 = _GEN_11958 & _GEN_12025 ? 1'h0 : _GEN_3373; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4406 = _GEN_11958 & _GEN_12027 ? 1'h0 : _GEN_3374; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4407 = _GEN_11958 & _GEN_12029 ? 1'h0 : _GEN_3375; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4408 = _GEN_11958 & _GEN_12031 ? 1'h0 : _GEN_3376; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4409 = _GEN_11958 & _GEN_12033 ? 1'h0 : _GEN_3377; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4410 = _GEN_11958 & _GEN_12035 ? 1'h0 : _GEN_3378; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4411 = _GEN_11958 & _GEN_12037 ? 1'h0 : _GEN_3379; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4412 = _GEN_11958 & _GEN_12039 ? 1'h0 : _GEN_3380; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4413 = _GEN_11958 & _GEN_12041 ? 1'h0 : _GEN_3381; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4414 = _GEN_11958 & _GEN_12043 ? 1'h0 : _GEN_3382; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4415 = _GEN_11958 & _GEN_12045 ? 1'h0 : _GEN_3383; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4416 = _GEN_11958 & _GEN_12047 ? 1'h0 : _GEN_3384; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4417 = _GEN_11958 & _GEN_12049 ? 1'h0 : _GEN_3385; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4418 = _GEN_11958 & _GEN_12051 ? 1'h0 : _GEN_3386; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4419 = _GEN_11958 & _GEN_12053 ? 1'h0 : _GEN_3387; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4420 = _GEN_11958 & _GEN_12055 ? 1'h0 : _GEN_3388; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4421 = _GEN_11958 & _GEN_12057 ? 1'h0 : _GEN_3389; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4422 = _GEN_11958 & _GEN_12059 ? 1'h0 : _GEN_3390; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4423 = _GEN_11958 & _GEN_12061 ? 1'h0 : _GEN_3391; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4424 = _GEN_11958 & _GEN_12063 ? 1'h0 : _GEN_3392; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4425 = _GEN_11958 & _GEN_12065 ? 1'h0 : _GEN_3393; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4426 = _GEN_11958 & _GEN_12067 ? 1'h0 : _GEN_3394; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4427 = _GEN_11958 & _GEN_12069 ? 1'h0 : _GEN_3395; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4428 = _GEN_11958 & _GEN_12071 ? 1'h0 : _GEN_3396; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4429 = _GEN_11958 & _GEN_12073 ? 1'h0 : _GEN_3397; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4430 = _GEN_11958 & _GEN_12075 ? 1'h0 : _GEN_3398; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4431 = _GEN_11958 & _GEN_12077 ? 1'h0 : _GEN_3399; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4432 = _GEN_11958 & _GEN_12079 ? 1'h0 : _GEN_3400; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4433 = _GEN_11958 & _GEN_12081 ? 1'h0 : _GEN_3401; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4434 = _GEN_11958 & _GEN_12083 ? 1'h0 : _GEN_3402; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4435 = _GEN_11958 & _GEN_12085 ? 1'h0 : _GEN_3403; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4436 = _GEN_11958 & _GEN_12087 ? 1'h0 : _GEN_3404; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4437 = _GEN_11958 & _GEN_12089 ? 1'h0 : _GEN_3405; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4438 = _GEN_11958 & _GEN_12091 ? 1'h0 : _GEN_3406; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4439 = _GEN_11958 & _GEN_12093 ? 1'h0 : _GEN_3407; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4440 = _GEN_11958 & _GEN_12095 ? 1'h0 : _GEN_3408; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4441 = _GEN_11958 & _GEN_12097 ? 1'h0 : _GEN_3409; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4442 = _GEN_11958 & _GEN_12099 ? 1'h0 : _GEN_3410; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4443 = _GEN_11958 & _GEN_12101 ? 1'h0 : _GEN_3411; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4444 = _GEN_11958 & _GEN_12103 ? 1'h0 : _GEN_3412; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4445 = _GEN_11958 & _GEN_12105 ? 1'h0 : _GEN_3413; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4446 = _GEN_11958 & _GEN_12107 ? 1'h0 : _GEN_3414; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4447 = _GEN_11958 & _GEN_12109 ? 1'h0 : _GEN_3415; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4448 = _GEN_11958 & _GEN_12111 ? 1'h0 : _GEN_3416; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4449 = _GEN_11958 & _GEN_12113 ? 1'h0 : _GEN_3417; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4450 = _GEN_11958 & _GEN_12115 ? 1'h0 : _GEN_3418; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4451 = _GEN_11958 & _GEN_12117 ? 1'h0 : _GEN_3419; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4452 = _GEN_11958 & _GEN_12119 ? 1'h0 : _GEN_3420; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4453 = _GEN_11958 & _GEN_12121 ? 1'h0 : _GEN_3421; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4454 = _GEN_11958 & _GEN_12123 ? 1'h0 : _GEN_3422; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4455 = _GEN_11958 & _GEN_12125 ? 1'h0 : _GEN_3423; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4456 = _GEN_11958 & _GEN_12127 ? 1'h0 : _GEN_3424; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4457 = _GEN_11958 & _GEN_12129 ? 1'h0 : _GEN_3425; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4458 = _GEN_11958 & _GEN_12131 ? 1'h0 : _GEN_3426; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4459 = _GEN_11958 & _GEN_12133 ? 1'h0 : _GEN_3427; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4460 = _GEN_11958 & _GEN_12135 ? 1'h0 : _GEN_3428; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4461 = _GEN_11958 & _GEN_12137 ? 1'h0 : _GEN_3429; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4462 = _GEN_11958 & _GEN_12139 ? 1'h0 : _GEN_3430; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4463 = _GEN_11958 & _GEN_12141 ? 1'h0 : _GEN_3431; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4464 = _GEN_11958 & _GEN_12143 ? 1'h0 : _GEN_3432; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4465 = _GEN_11958 & _GEN_12145 ? 1'h0 : _GEN_3433; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4466 = _GEN_11958 & _GEN_12147 ? 1'h0 : _GEN_3434; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4467 = _GEN_11958 & _GEN_12149 ? 1'h0 : _GEN_3435; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4468 = _GEN_11958 & _GEN_12151 ? 1'h0 : _GEN_3436; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4469 = _GEN_11958 & _GEN_12153 ? 1'h0 : _GEN_3437; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4470 = _GEN_11958 & _GEN_12155 ? 1'h0 : _GEN_3438; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4471 = _GEN_11958 & _GEN_12157 ? 1'h0 : _GEN_3439; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4472 = _GEN_11958 & _GEN_12159 ? 1'h0 : _GEN_3440; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4473 = _GEN_11958 & _GEN_12161 ? 1'h0 : _GEN_3441; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4474 = _GEN_11958 & _GEN_12163 ? 1'h0 : _GEN_3442; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4475 = _GEN_11958 & _GEN_12165 ? 1'h0 : _GEN_3443; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4476 = _GEN_11958 & _GEN_12167 ? 1'h0 : _GEN_3444; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4477 = _GEN_11958 & _GEN_12169 ? 1'h0 : _GEN_3445; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4478 = _GEN_11958 & _GEN_12171 ? 1'h0 : _GEN_3446; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4479 = _GEN_11958 & _GEN_12173 ? 1'h0 : _GEN_3447; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4480 = _GEN_11958 & _GEN_12175 ? 1'h0 : _GEN_3448; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4481 = _GEN_11958 & _GEN_12177 ? 1'h0 : _GEN_3449; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4482 = _GEN_11958 & _GEN_12179 ? 1'h0 : _GEN_3450; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4483 = _GEN_11958 & _GEN_12181 ? 1'h0 : _GEN_3451; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4484 = _GEN_11958 & _GEN_12183 ? 1'h0 : _GEN_3452; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4485 = _GEN_11958 & _GEN_12185 ? 1'h0 : _GEN_3453; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4486 = _GEN_11958 & _GEN_12187 ? 1'h0 : _GEN_3454; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4487 = _GEN_11958 & _GEN_12189 ? 1'h0 : _GEN_3455; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4488 = _GEN_11958 & _GEN_12191 ? 1'h0 : _GEN_3456; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4489 = _GEN_11958 & _GEN_12193 ? 1'h0 : _GEN_3457; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4490 = _GEN_11958 & _GEN_12195 ? 1'h0 : _GEN_3458; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4491 = _GEN_11958 & _GEN_12197 ? 1'h0 : _GEN_3459; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4492 = _GEN_11958 & _GEN_12199 ? 1'h0 : _GEN_3460; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4493 = _GEN_11958 & _GEN_12201 ? 1'h0 : _GEN_3461; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4494 = _GEN_11958 & _GEN_12203 ? 1'h0 : _GEN_3462; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4495 = _GEN_11958 & _GEN_12205 ? 1'h0 : _GEN_3463; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4496 = _GEN_11958 & _GEN_12207 ? 1'h0 : _GEN_3464; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4497 = _GEN_11958 & _GEN_12209 ? 1'h0 : _GEN_3465; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4498 = _GEN_11958 & _GEN_12211 ? 1'h0 : _GEN_3466; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4499 = _GEN_11958 & _GEN_12213 ? 1'h0 : _GEN_3467; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4500 = _GEN_11958 & _GEN_12215 ? 1'h0 : _GEN_3468; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4501 = _GEN_11958 & _GEN_12217 ? 1'h0 : _GEN_3469; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4502 = _GEN_11958 & _GEN_12219 ? 1'h0 : _GEN_3470; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4503 = _GEN_11958 & _GEN_12221 ? 1'h0 : _GEN_3471; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4504 = _GEN_11958 & _GEN_12223 ? 1'h0 : _GEN_3472; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4505 = _GEN_11958 & _GEN_12225 ? 1'h0 : _GEN_3473; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4506 = _GEN_11958 & _GEN_12227 ? 1'h0 : _GEN_3474; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4507 = _GEN_11958 & _GEN_12229 ? 1'h0 : _GEN_3475; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4508 = _GEN_11958 & _GEN_12231 ? 1'h0 : _GEN_3476; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4509 = _GEN_11958 & _GEN_12233 ? 1'h0 : _GEN_3477; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4510 = _GEN_11958 & _GEN_12235 ? 1'h0 : _GEN_3478; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4511 = _GEN_11958 & _GEN_12237 ? 1'h0 : _GEN_3479; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4512 = _GEN_11958 & _GEN_12239 ? 1'h0 : _GEN_3480; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4513 = _GEN_11958 & _GEN_12241 ? 1'h0 : _GEN_3481; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4514 = _GEN_11958 & _GEN_12243 ? 1'h0 : _GEN_3482; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4515 = _GEN_11958 & _GEN_12245 ? 1'h0 : _GEN_3483; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4516 = _GEN_11958 & _GEN_12247 ? 1'h0 : _GEN_3484; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4517 = _GEN_11958 & _GEN_12249 ? 1'h0 : _GEN_3485; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4518 = _GEN_11958 & _GEN_12251 ? 1'h0 : _GEN_3486; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4519 = _GEN_11958 & _GEN_12253 ? 1'h0 : _GEN_3487; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4520 = _GEN_11958 & _GEN_12255 ? 1'h0 : _GEN_3488; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4521 = _GEN_11958 & _GEN_12257 ? 1'h0 : _GEN_3489; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4522 = _GEN_11958 & _GEN_12259 ? 1'h0 : _GEN_3490; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4523 = _GEN_11958 & _GEN_12261 ? 1'h0 : _GEN_3491; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4524 = _GEN_11958 & _GEN_12263 ? 1'h0 : _GEN_3492; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4525 = _GEN_11958 & _GEN_12265 ? 1'h0 : _GEN_3493; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4526 = _GEN_11958 & _GEN_12267 ? 1'h0 : _GEN_3494; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4527 = _GEN_11958 & _GEN_12269 ? 1'h0 : _GEN_3495; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4528 = _GEN_11958 & _GEN_12271 ? 1'h0 : _GEN_3496; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4529 = _GEN_11958 & _GEN_12273 ? 1'h0 : _GEN_3497; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4530 = _GEN_11958 & _GEN_12275 ? 1'h0 : _GEN_3498; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4531 = _GEN_11958 & _GEN_12277 ? 1'h0 : _GEN_3499; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4532 = _GEN_11958 & _GEN_12279 ? 1'h0 : _GEN_3500; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4533 = _GEN_11958 & _GEN_12281 ? 1'h0 : _GEN_3501; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4534 = _GEN_11958 & _GEN_12283 ? 1'h0 : _GEN_3502; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4535 = _GEN_11958 & _GEN_12285 ? 1'h0 : _GEN_3503; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4536 = _GEN_11958 & _GEN_12287 ? 1'h0 : _GEN_3504; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4537 = _GEN_11958 & _GEN_12289 ? 1'h0 : _GEN_3505; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4538 = _GEN_11958 & _GEN_12291 ? 1'h0 : _GEN_3506; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4539 = _GEN_11958 & _GEN_12293 ? 1'h0 : _GEN_3507; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4540 = _GEN_11958 & _GEN_12295 ? 1'h0 : _GEN_3508; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4541 = _GEN_11958 & _GEN_12297 ? 1'h0 : _GEN_3509; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4542 = _GEN_11958 & _GEN_12299 ? 1'h0 : _GEN_3510; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4543 = _GEN_11958 & _GEN_12301 ? 1'h0 : _GEN_3511; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4544 = _GEN_11958 & _GEN_12303 ? 1'h0 : _GEN_3512; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4545 = _GEN_11958 & _GEN_12305 ? 1'h0 : _GEN_3513; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4546 = _GEN_11958 & _GEN_12307 ? 1'h0 : _GEN_3514; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4547 = _GEN_11958 & _GEN_12309 ? 1'h0 : _GEN_3515; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4548 = _GEN_11958 & _GEN_12311 ? 1'h0 : _GEN_3516; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4549 = _GEN_11958 & _GEN_12313 ? 1'h0 : _GEN_3517; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4550 = _GEN_11958 & _GEN_12315 ? 1'h0 : _GEN_3518; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4551 = _GEN_11958 & _GEN_12317 ? 1'h0 : _GEN_3519; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4552 = _GEN_11958 & _GEN_12319 ? 1'h0 : _GEN_3520; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4553 = _GEN_11958 & _GEN_12321 ? 1'h0 : _GEN_3521; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4554 = _GEN_11958 & _GEN_12323 ? 1'h0 : _GEN_3522; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4555 = _GEN_11958 & _GEN_12325 ? 1'h0 : _GEN_3523; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4556 = _GEN_11958 & _GEN_12327 ? 1'h0 : _GEN_3524; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4557 = _GEN_11958 & _GEN_12329 ? 1'h0 : _GEN_3525; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4558 = _GEN_11958 & _GEN_12331 ? 1'h0 : _GEN_3526; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4559 = _GEN_11958 & _GEN_12333 ? 1'h0 : _GEN_3527; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4560 = _GEN_11958 & _GEN_12335 ? 1'h0 : _GEN_3528; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4561 = _GEN_11958 & _GEN_12337 ? 1'h0 : _GEN_3529; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4562 = _GEN_11958 & _GEN_12339 ? 1'h0 : _GEN_3530; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4563 = _GEN_11958 & _GEN_12341 ? 1'h0 : _GEN_3531; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4564 = _GEN_11958 & _GEN_12343 ? 1'h0 : _GEN_3532; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4565 = _GEN_11958 & _GEN_12345 ? 1'h0 : _GEN_3533; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4566 = _GEN_11958 & _GEN_12347 ? 1'h0 : _GEN_3534; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4567 = _GEN_11958 & _GEN_12349 ? 1'h0 : _GEN_3535; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4568 = _GEN_11958 & _GEN_12351 ? 1'h0 : _GEN_3536; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4569 = _GEN_11958 & _GEN_12353 ? 1'h0 : _GEN_3537; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4570 = _GEN_11958 & _GEN_12355 ? 1'h0 : _GEN_3538; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4571 = _GEN_11958 & _GEN_12357 ? 1'h0 : _GEN_3539; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4572 = _GEN_11958 & _GEN_12359 ? 1'h0 : _GEN_3540; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4573 = _GEN_11958 & _GEN_12361 ? 1'h0 : _GEN_3541; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4574 = _GEN_11958 & _GEN_12363 ? 1'h0 : _GEN_3542; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4575 = _GEN_11958 & _GEN_12365 ? 1'h0 : _GEN_3543; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4576 = _GEN_11958 & _GEN_12367 ? 1'h0 : _GEN_3544; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4577 = _GEN_11958 & _GEN_12369 ? 1'h0 : _GEN_3545; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4578 = _GEN_11958 & _GEN_12371 ? 1'h0 : _GEN_3546; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4579 = _GEN_11958 & _GEN_12373 ? 1'h0 : _GEN_3547; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4580 = _GEN_11958 & _GEN_12375 ? 1'h0 : _GEN_3548; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4581 = _GEN_11958 & _GEN_12377 ? 1'h0 : _GEN_3549; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4582 = _GEN_11958 & _GEN_12379 ? 1'h0 : _GEN_3550; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4583 = _GEN_11958 & _GEN_12381 ? 1'h0 : _GEN_3551; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4584 = _GEN_11958 & _GEN_12383 ? 1'h0 : _GEN_3552; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4585 = _GEN_11958 & _GEN_12385 ? 1'h0 : _GEN_3553; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4586 = _GEN_11958 & _GEN_12387 ? 1'h0 : _GEN_3554; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4587 = _GEN_11958 & _GEN_12389 ? 1'h0 : _GEN_3555; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4588 = _GEN_11958 & _GEN_12391 ? 1'h0 : _GEN_3556; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4589 = _GEN_11958 & _GEN_12393 ? 1'h0 : _GEN_3557; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4590 = _GEN_11958 & _GEN_12395 ? 1'h0 : _GEN_3558; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4591 = _GEN_11958 & _GEN_12397 ? 1'h0 : _GEN_3559; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4592 = _GEN_11958 & _GEN_12399 ? 1'h0 : _GEN_3560; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4593 = _GEN_11958 & _GEN_12401 ? 1'h0 : _GEN_3561; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4594 = _GEN_11958 & _GEN_12403 ? 1'h0 : _GEN_3562; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4595 = _GEN_11958 & _GEN_12405 ? 1'h0 : _GEN_3563; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4596 = _GEN_11958 & _GEN_12407 ? 1'h0 : _GEN_3564; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4597 = _GEN_11958 & _GEN_12409 ? 1'h0 : _GEN_3565; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4598 = _GEN_11958 & _GEN_12411 ? 1'h0 : _GEN_3566; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4599 = _GEN_11958 & _GEN_12413 ? 1'h0 : _GEN_3567; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4600 = _GEN_11958 & _GEN_12415 ? 1'h0 : _GEN_3568; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4601 = _GEN_11958 & _GEN_12417 ? 1'h0 : _GEN_3569; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4602 = _GEN_11958 & _GEN_12419 ? 1'h0 : _GEN_3570; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4603 = _GEN_11958 & _GEN_12421 ? 1'h0 : _GEN_3571; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4604 = _GEN_11958 & _GEN_12423 ? 1'h0 : _GEN_3572; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4605 = _GEN_11958 & _GEN_12425 ? 1'h0 : _GEN_3573; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4606 = _GEN_11958 & _GEN_12427 ? 1'h0 : _GEN_3574; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4607 = _GEN_11958 & _GEN_12429 ? 1'h0 : _GEN_3575; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4608 = _GEN_11958 & _GEN_12431 ? 1'h0 : _GEN_3576; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4609 = _GEN_11958 & _GEN_12433 ? 1'h0 : _GEN_3577; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4610 = _GEN_11958 & _GEN_12435 ? 1'h0 : _GEN_3578; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4611 = _GEN_11958 & _GEN_12437 ? 1'h0 : _GEN_3579; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4612 = _GEN_11958 & _GEN_12439 ? 1'h0 : _GEN_3580; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4613 = _GEN_11958 & _GEN_12441 ? 1'h0 : _GEN_3581; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4614 = _GEN_11958 & _GEN_12443 ? 1'h0 : _GEN_3582; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4615 = _GEN_11958 & _GEN_12445 ? 1'h0 : _GEN_3583; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4616 = _GEN_11958 & _GEN_12447 ? 1'h0 : _GEN_3584; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4617 = _GEN_11958 & _GEN_12449 ? 1'h0 : _GEN_3585; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4618 = _GEN_11958 & _GEN_12451 ? 1'h0 : _GEN_3586; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4619 = _GEN_11958 & _GEN_12453 ? 1'h0 : _GEN_3587; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4620 = _GEN_11958 & _GEN_12455 ? 1'h0 : _GEN_3588; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4621 = _GEN_11958 & _GEN_12457 ? 1'h0 : _GEN_3589; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4622 = _GEN_11958 & _GEN_12459 ? 1'h0 : _GEN_3590; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4623 = _GEN_11958 & _GEN_12461 ? 1'h0 : _GEN_3591; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4624 = _GEN_11958 & _GEN_12463 ? 1'h0 : _GEN_3592; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4625 = _GEN_11958 & _GEN_12465 ? 1'h0 : _GEN_3593; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4626 = _GEN_11958 & _GEN_12467 ? 1'h0 : _GEN_3594; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4627 = refillIDX_r & _GEN_12468 ? 1'h0 : _GEN_3595; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4628 = refillIDX_r & _GEN_11959 ? 1'h0 : _GEN_3596; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4629 = refillIDX_r & _GEN_11961 ? 1'h0 : _GEN_3597; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4630 = refillIDX_r & _GEN_11963 ? 1'h0 : _GEN_3598; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4631 = refillIDX_r & _GEN_11965 ? 1'h0 : _GEN_3599; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4632 = refillIDX_r & _GEN_11967 ? 1'h0 : _GEN_3600; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4633 = refillIDX_r & _GEN_11969 ? 1'h0 : _GEN_3601; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4634 = refillIDX_r & _GEN_11971 ? 1'h0 : _GEN_3602; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4635 = refillIDX_r & _GEN_11973 ? 1'h0 : _GEN_3603; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4636 = refillIDX_r & _GEN_11975 ? 1'h0 : _GEN_3604; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4637 = refillIDX_r & _GEN_11977 ? 1'h0 : _GEN_3605; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4638 = refillIDX_r & _GEN_11979 ? 1'h0 : _GEN_3606; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4639 = refillIDX_r & _GEN_11981 ? 1'h0 : _GEN_3607; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4640 = refillIDX_r & _GEN_11983 ? 1'h0 : _GEN_3608; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4641 = refillIDX_r & _GEN_11985 ? 1'h0 : _GEN_3609; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4642 = refillIDX_r & _GEN_11987 ? 1'h0 : _GEN_3610; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4643 = refillIDX_r & _GEN_11989 ? 1'h0 : _GEN_3611; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4644 = refillIDX_r & _GEN_11991 ? 1'h0 : _GEN_3612; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4645 = refillIDX_r & _GEN_11993 ? 1'h0 : _GEN_3613; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4646 = refillIDX_r & _GEN_11995 ? 1'h0 : _GEN_3614; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4647 = refillIDX_r & _GEN_11997 ? 1'h0 : _GEN_3615; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4648 = refillIDX_r & _GEN_11999 ? 1'h0 : _GEN_3616; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4649 = refillIDX_r & _GEN_12001 ? 1'h0 : _GEN_3617; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4650 = refillIDX_r & _GEN_12003 ? 1'h0 : _GEN_3618; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4651 = refillIDX_r & _GEN_12005 ? 1'h0 : _GEN_3619; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4652 = refillIDX_r & _GEN_12007 ? 1'h0 : _GEN_3620; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4653 = refillIDX_r & _GEN_12009 ? 1'h0 : _GEN_3621; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4654 = refillIDX_r & _GEN_12011 ? 1'h0 : _GEN_3622; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4655 = refillIDX_r & _GEN_12013 ? 1'h0 : _GEN_3623; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4656 = refillIDX_r & _GEN_12015 ? 1'h0 : _GEN_3624; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4657 = refillIDX_r & _GEN_12017 ? 1'h0 : _GEN_3625; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4658 = refillIDX_r & _GEN_12019 ? 1'h0 : _GEN_3626; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4659 = refillIDX_r & _GEN_12021 ? 1'h0 : _GEN_3627; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4660 = refillIDX_r & _GEN_12023 ? 1'h0 : _GEN_3628; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4661 = refillIDX_r & _GEN_12025 ? 1'h0 : _GEN_3629; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4662 = refillIDX_r & _GEN_12027 ? 1'h0 : _GEN_3630; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4663 = refillIDX_r & _GEN_12029 ? 1'h0 : _GEN_3631; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4664 = refillIDX_r & _GEN_12031 ? 1'h0 : _GEN_3632; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4665 = refillIDX_r & _GEN_12033 ? 1'h0 : _GEN_3633; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4666 = refillIDX_r & _GEN_12035 ? 1'h0 : _GEN_3634; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4667 = refillIDX_r & _GEN_12037 ? 1'h0 : _GEN_3635; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4668 = refillIDX_r & _GEN_12039 ? 1'h0 : _GEN_3636; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4669 = refillIDX_r & _GEN_12041 ? 1'h0 : _GEN_3637; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4670 = refillIDX_r & _GEN_12043 ? 1'h0 : _GEN_3638; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4671 = refillIDX_r & _GEN_12045 ? 1'h0 : _GEN_3639; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4672 = refillIDX_r & _GEN_12047 ? 1'h0 : _GEN_3640; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4673 = refillIDX_r & _GEN_12049 ? 1'h0 : _GEN_3641; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4674 = refillIDX_r & _GEN_12051 ? 1'h0 : _GEN_3642; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4675 = refillIDX_r & _GEN_12053 ? 1'h0 : _GEN_3643; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4676 = refillIDX_r & _GEN_12055 ? 1'h0 : _GEN_3644; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4677 = refillIDX_r & _GEN_12057 ? 1'h0 : _GEN_3645; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4678 = refillIDX_r & _GEN_12059 ? 1'h0 : _GEN_3646; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4679 = refillIDX_r & _GEN_12061 ? 1'h0 : _GEN_3647; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4680 = refillIDX_r & _GEN_12063 ? 1'h0 : _GEN_3648; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4681 = refillIDX_r & _GEN_12065 ? 1'h0 : _GEN_3649; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4682 = refillIDX_r & _GEN_12067 ? 1'h0 : _GEN_3650; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4683 = refillIDX_r & _GEN_12069 ? 1'h0 : _GEN_3651; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4684 = refillIDX_r & _GEN_12071 ? 1'h0 : _GEN_3652; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4685 = refillIDX_r & _GEN_12073 ? 1'h0 : _GEN_3653; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4686 = refillIDX_r & _GEN_12075 ? 1'h0 : _GEN_3654; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4687 = refillIDX_r & _GEN_12077 ? 1'h0 : _GEN_3655; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4688 = refillIDX_r & _GEN_12079 ? 1'h0 : _GEN_3656; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4689 = refillIDX_r & _GEN_12081 ? 1'h0 : _GEN_3657; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4690 = refillIDX_r & _GEN_12083 ? 1'h0 : _GEN_3658; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4691 = refillIDX_r & _GEN_12085 ? 1'h0 : _GEN_3659; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4692 = refillIDX_r & _GEN_12087 ? 1'h0 : _GEN_3660; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4693 = refillIDX_r & _GEN_12089 ? 1'h0 : _GEN_3661; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4694 = refillIDX_r & _GEN_12091 ? 1'h0 : _GEN_3662; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4695 = refillIDX_r & _GEN_12093 ? 1'h0 : _GEN_3663; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4696 = refillIDX_r & _GEN_12095 ? 1'h0 : _GEN_3664; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4697 = refillIDX_r & _GEN_12097 ? 1'h0 : _GEN_3665; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4698 = refillIDX_r & _GEN_12099 ? 1'h0 : _GEN_3666; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4699 = refillIDX_r & _GEN_12101 ? 1'h0 : _GEN_3667; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4700 = refillIDX_r & _GEN_12103 ? 1'h0 : _GEN_3668; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4701 = refillIDX_r & _GEN_12105 ? 1'h0 : _GEN_3669; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4702 = refillIDX_r & _GEN_12107 ? 1'h0 : _GEN_3670; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4703 = refillIDX_r & _GEN_12109 ? 1'h0 : _GEN_3671; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4704 = refillIDX_r & _GEN_12111 ? 1'h0 : _GEN_3672; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4705 = refillIDX_r & _GEN_12113 ? 1'h0 : _GEN_3673; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4706 = refillIDX_r & _GEN_12115 ? 1'h0 : _GEN_3674; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4707 = refillIDX_r & _GEN_12117 ? 1'h0 : _GEN_3675; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4708 = refillIDX_r & _GEN_12119 ? 1'h0 : _GEN_3676; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4709 = refillIDX_r & _GEN_12121 ? 1'h0 : _GEN_3677; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4710 = refillIDX_r & _GEN_12123 ? 1'h0 : _GEN_3678; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4711 = refillIDX_r & _GEN_12125 ? 1'h0 : _GEN_3679; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4712 = refillIDX_r & _GEN_12127 ? 1'h0 : _GEN_3680; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4713 = refillIDX_r & _GEN_12129 ? 1'h0 : _GEN_3681; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4714 = refillIDX_r & _GEN_12131 ? 1'h0 : _GEN_3682; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4715 = refillIDX_r & _GEN_12133 ? 1'h0 : _GEN_3683; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4716 = refillIDX_r & _GEN_12135 ? 1'h0 : _GEN_3684; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4717 = refillIDX_r & _GEN_12137 ? 1'h0 : _GEN_3685; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4718 = refillIDX_r & _GEN_12139 ? 1'h0 : _GEN_3686; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4719 = refillIDX_r & _GEN_12141 ? 1'h0 : _GEN_3687; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4720 = refillIDX_r & _GEN_12143 ? 1'h0 : _GEN_3688; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4721 = refillIDX_r & _GEN_12145 ? 1'h0 : _GEN_3689; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4722 = refillIDX_r & _GEN_12147 ? 1'h0 : _GEN_3690; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4723 = refillIDX_r & _GEN_12149 ? 1'h0 : _GEN_3691; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4724 = refillIDX_r & _GEN_12151 ? 1'h0 : _GEN_3692; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4725 = refillIDX_r & _GEN_12153 ? 1'h0 : _GEN_3693; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4726 = refillIDX_r & _GEN_12155 ? 1'h0 : _GEN_3694; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4727 = refillIDX_r & _GEN_12157 ? 1'h0 : _GEN_3695; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4728 = refillIDX_r & _GEN_12159 ? 1'h0 : _GEN_3696; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4729 = refillIDX_r & _GEN_12161 ? 1'h0 : _GEN_3697; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4730 = refillIDX_r & _GEN_12163 ? 1'h0 : _GEN_3698; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4731 = refillIDX_r & _GEN_12165 ? 1'h0 : _GEN_3699; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4732 = refillIDX_r & _GEN_12167 ? 1'h0 : _GEN_3700; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4733 = refillIDX_r & _GEN_12169 ? 1'h0 : _GEN_3701; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4734 = refillIDX_r & _GEN_12171 ? 1'h0 : _GEN_3702; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4735 = refillIDX_r & _GEN_12173 ? 1'h0 : _GEN_3703; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4736 = refillIDX_r & _GEN_12175 ? 1'h0 : _GEN_3704; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4737 = refillIDX_r & _GEN_12177 ? 1'h0 : _GEN_3705; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4738 = refillIDX_r & _GEN_12179 ? 1'h0 : _GEN_3706; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4739 = refillIDX_r & _GEN_12181 ? 1'h0 : _GEN_3707; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4740 = refillIDX_r & _GEN_12183 ? 1'h0 : _GEN_3708; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4741 = refillIDX_r & _GEN_12185 ? 1'h0 : _GEN_3709; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4742 = refillIDX_r & _GEN_12187 ? 1'h0 : _GEN_3710; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4743 = refillIDX_r & _GEN_12189 ? 1'h0 : _GEN_3711; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4744 = refillIDX_r & _GEN_12191 ? 1'h0 : _GEN_3712; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4745 = refillIDX_r & _GEN_12193 ? 1'h0 : _GEN_3713; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4746 = refillIDX_r & _GEN_12195 ? 1'h0 : _GEN_3714; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4747 = refillIDX_r & _GEN_12197 ? 1'h0 : _GEN_3715; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4748 = refillIDX_r & _GEN_12199 ? 1'h0 : _GEN_3716; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4749 = refillIDX_r & _GEN_12201 ? 1'h0 : _GEN_3717; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4750 = refillIDX_r & _GEN_12203 ? 1'h0 : _GEN_3718; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4751 = refillIDX_r & _GEN_12205 ? 1'h0 : _GEN_3719; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4752 = refillIDX_r & _GEN_12207 ? 1'h0 : _GEN_3720; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4753 = refillIDX_r & _GEN_12209 ? 1'h0 : _GEN_3721; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4754 = refillIDX_r & _GEN_12211 ? 1'h0 : _GEN_3722; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4755 = refillIDX_r & _GEN_12213 ? 1'h0 : _GEN_3723; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4756 = refillIDX_r & _GEN_12215 ? 1'h0 : _GEN_3724; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4757 = refillIDX_r & _GEN_12217 ? 1'h0 : _GEN_3725; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4758 = refillIDX_r & _GEN_12219 ? 1'h0 : _GEN_3726; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4759 = refillIDX_r & _GEN_12221 ? 1'h0 : _GEN_3727; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4760 = refillIDX_r & _GEN_12223 ? 1'h0 : _GEN_3728; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4761 = refillIDX_r & _GEN_12225 ? 1'h0 : _GEN_3729; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4762 = refillIDX_r & _GEN_12227 ? 1'h0 : _GEN_3730; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4763 = refillIDX_r & _GEN_12229 ? 1'h0 : _GEN_3731; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4764 = refillIDX_r & _GEN_12231 ? 1'h0 : _GEN_3732; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4765 = refillIDX_r & _GEN_12233 ? 1'h0 : _GEN_3733; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4766 = refillIDX_r & _GEN_12235 ? 1'h0 : _GEN_3734; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4767 = refillIDX_r & _GEN_12237 ? 1'h0 : _GEN_3735; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4768 = refillIDX_r & _GEN_12239 ? 1'h0 : _GEN_3736; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4769 = refillIDX_r & _GEN_12241 ? 1'h0 : _GEN_3737; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4770 = refillIDX_r & _GEN_12243 ? 1'h0 : _GEN_3738; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4771 = refillIDX_r & _GEN_12245 ? 1'h0 : _GEN_3739; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4772 = refillIDX_r & _GEN_12247 ? 1'h0 : _GEN_3740; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4773 = refillIDX_r & _GEN_12249 ? 1'h0 : _GEN_3741; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4774 = refillIDX_r & _GEN_12251 ? 1'h0 : _GEN_3742; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4775 = refillIDX_r & _GEN_12253 ? 1'h0 : _GEN_3743; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4776 = refillIDX_r & _GEN_12255 ? 1'h0 : _GEN_3744; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4777 = refillIDX_r & _GEN_12257 ? 1'h0 : _GEN_3745; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4778 = refillIDX_r & _GEN_12259 ? 1'h0 : _GEN_3746; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4779 = refillIDX_r & _GEN_12261 ? 1'h0 : _GEN_3747; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4780 = refillIDX_r & _GEN_12263 ? 1'h0 : _GEN_3748; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4781 = refillIDX_r & _GEN_12265 ? 1'h0 : _GEN_3749; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4782 = refillIDX_r & _GEN_12267 ? 1'h0 : _GEN_3750; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4783 = refillIDX_r & _GEN_12269 ? 1'h0 : _GEN_3751; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4784 = refillIDX_r & _GEN_12271 ? 1'h0 : _GEN_3752; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4785 = refillIDX_r & _GEN_12273 ? 1'h0 : _GEN_3753; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4786 = refillIDX_r & _GEN_12275 ? 1'h0 : _GEN_3754; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4787 = refillIDX_r & _GEN_12277 ? 1'h0 : _GEN_3755; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4788 = refillIDX_r & _GEN_12279 ? 1'h0 : _GEN_3756; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4789 = refillIDX_r & _GEN_12281 ? 1'h0 : _GEN_3757; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4790 = refillIDX_r & _GEN_12283 ? 1'h0 : _GEN_3758; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4791 = refillIDX_r & _GEN_12285 ? 1'h0 : _GEN_3759; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4792 = refillIDX_r & _GEN_12287 ? 1'h0 : _GEN_3760; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4793 = refillIDX_r & _GEN_12289 ? 1'h0 : _GEN_3761; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4794 = refillIDX_r & _GEN_12291 ? 1'h0 : _GEN_3762; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4795 = refillIDX_r & _GEN_12293 ? 1'h0 : _GEN_3763; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4796 = refillIDX_r & _GEN_12295 ? 1'h0 : _GEN_3764; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4797 = refillIDX_r & _GEN_12297 ? 1'h0 : _GEN_3765; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4798 = refillIDX_r & _GEN_12299 ? 1'h0 : _GEN_3766; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4799 = refillIDX_r & _GEN_12301 ? 1'h0 : _GEN_3767; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4800 = refillIDX_r & _GEN_12303 ? 1'h0 : _GEN_3768; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4801 = refillIDX_r & _GEN_12305 ? 1'h0 : _GEN_3769; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4802 = refillIDX_r & _GEN_12307 ? 1'h0 : _GEN_3770; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4803 = refillIDX_r & _GEN_12309 ? 1'h0 : _GEN_3771; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4804 = refillIDX_r & _GEN_12311 ? 1'h0 : _GEN_3772; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4805 = refillIDX_r & _GEN_12313 ? 1'h0 : _GEN_3773; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4806 = refillIDX_r & _GEN_12315 ? 1'h0 : _GEN_3774; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4807 = refillIDX_r & _GEN_12317 ? 1'h0 : _GEN_3775; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4808 = refillIDX_r & _GEN_12319 ? 1'h0 : _GEN_3776; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4809 = refillIDX_r & _GEN_12321 ? 1'h0 : _GEN_3777; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4810 = refillIDX_r & _GEN_12323 ? 1'h0 : _GEN_3778; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4811 = refillIDX_r & _GEN_12325 ? 1'h0 : _GEN_3779; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4812 = refillIDX_r & _GEN_12327 ? 1'h0 : _GEN_3780; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4813 = refillIDX_r & _GEN_12329 ? 1'h0 : _GEN_3781; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4814 = refillIDX_r & _GEN_12331 ? 1'h0 : _GEN_3782; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4815 = refillIDX_r & _GEN_12333 ? 1'h0 : _GEN_3783; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4816 = refillIDX_r & _GEN_12335 ? 1'h0 : _GEN_3784; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4817 = refillIDX_r & _GEN_12337 ? 1'h0 : _GEN_3785; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4818 = refillIDX_r & _GEN_12339 ? 1'h0 : _GEN_3786; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4819 = refillIDX_r & _GEN_12341 ? 1'h0 : _GEN_3787; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4820 = refillIDX_r & _GEN_12343 ? 1'h0 : _GEN_3788; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4821 = refillIDX_r & _GEN_12345 ? 1'h0 : _GEN_3789; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4822 = refillIDX_r & _GEN_12347 ? 1'h0 : _GEN_3790; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4823 = refillIDX_r & _GEN_12349 ? 1'h0 : _GEN_3791; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4824 = refillIDX_r & _GEN_12351 ? 1'h0 : _GEN_3792; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4825 = refillIDX_r & _GEN_12353 ? 1'h0 : _GEN_3793; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4826 = refillIDX_r & _GEN_12355 ? 1'h0 : _GEN_3794; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4827 = refillIDX_r & _GEN_12357 ? 1'h0 : _GEN_3795; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4828 = refillIDX_r & _GEN_12359 ? 1'h0 : _GEN_3796; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4829 = refillIDX_r & _GEN_12361 ? 1'h0 : _GEN_3797; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4830 = refillIDX_r & _GEN_12363 ? 1'h0 : _GEN_3798; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4831 = refillIDX_r & _GEN_12365 ? 1'h0 : _GEN_3799; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4832 = refillIDX_r & _GEN_12367 ? 1'h0 : _GEN_3800; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4833 = refillIDX_r & _GEN_12369 ? 1'h0 : _GEN_3801; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4834 = refillIDX_r & _GEN_12371 ? 1'h0 : _GEN_3802; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4835 = refillIDX_r & _GEN_12373 ? 1'h0 : _GEN_3803; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4836 = refillIDX_r & _GEN_12375 ? 1'h0 : _GEN_3804; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4837 = refillIDX_r & _GEN_12377 ? 1'h0 : _GEN_3805; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4838 = refillIDX_r & _GEN_12379 ? 1'h0 : _GEN_3806; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4839 = refillIDX_r & _GEN_12381 ? 1'h0 : _GEN_3807; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4840 = refillIDX_r & _GEN_12383 ? 1'h0 : _GEN_3808; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4841 = refillIDX_r & _GEN_12385 ? 1'h0 : _GEN_3809; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4842 = refillIDX_r & _GEN_12387 ? 1'h0 : _GEN_3810; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4843 = refillIDX_r & _GEN_12389 ? 1'h0 : _GEN_3811; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4844 = refillIDX_r & _GEN_12391 ? 1'h0 : _GEN_3812; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4845 = refillIDX_r & _GEN_12393 ? 1'h0 : _GEN_3813; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4846 = refillIDX_r & _GEN_12395 ? 1'h0 : _GEN_3814; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4847 = refillIDX_r & _GEN_12397 ? 1'h0 : _GEN_3815; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4848 = refillIDX_r & _GEN_12399 ? 1'h0 : _GEN_3816; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4849 = refillIDX_r & _GEN_12401 ? 1'h0 : _GEN_3817; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4850 = refillIDX_r & _GEN_12403 ? 1'h0 : _GEN_3818; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4851 = refillIDX_r & _GEN_12405 ? 1'h0 : _GEN_3819; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4852 = refillIDX_r & _GEN_12407 ? 1'h0 : _GEN_3820; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4853 = refillIDX_r & _GEN_12409 ? 1'h0 : _GEN_3821; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4854 = refillIDX_r & _GEN_12411 ? 1'h0 : _GEN_3822; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4855 = refillIDX_r & _GEN_12413 ? 1'h0 : _GEN_3823; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4856 = refillIDX_r & _GEN_12415 ? 1'h0 : _GEN_3824; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4857 = refillIDX_r & _GEN_12417 ? 1'h0 : _GEN_3825; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4858 = refillIDX_r & _GEN_12419 ? 1'h0 : _GEN_3826; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4859 = refillIDX_r & _GEN_12421 ? 1'h0 : _GEN_3827; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4860 = refillIDX_r & _GEN_12423 ? 1'h0 : _GEN_3828; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4861 = refillIDX_r & _GEN_12425 ? 1'h0 : _GEN_3829; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4862 = refillIDX_r & _GEN_12427 ? 1'h0 : _GEN_3830; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4863 = refillIDX_r & _GEN_12429 ? 1'h0 : _GEN_3831; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4864 = refillIDX_r & _GEN_12431 ? 1'h0 : _GEN_3832; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4865 = refillIDX_r & _GEN_12433 ? 1'h0 : _GEN_3833; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4866 = refillIDX_r & _GEN_12435 ? 1'h0 : _GEN_3834; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4867 = refillIDX_r & _GEN_12437 ? 1'h0 : _GEN_3835; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4868 = refillIDX_r & _GEN_12439 ? 1'h0 : _GEN_3836; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4869 = refillIDX_r & _GEN_12441 ? 1'h0 : _GEN_3837; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4870 = refillIDX_r & _GEN_12443 ? 1'h0 : _GEN_3838; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4871 = refillIDX_r & _GEN_12445 ? 1'h0 : _GEN_3839; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4872 = refillIDX_r & _GEN_12447 ? 1'h0 : _GEN_3840; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4873 = refillIDX_r & _GEN_12449 ? 1'h0 : _GEN_3841; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4874 = refillIDX_r & _GEN_12451 ? 1'h0 : _GEN_3842; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4875 = refillIDX_r & _GEN_12453 ? 1'h0 : _GEN_3843; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4876 = refillIDX_r & _GEN_12455 ? 1'h0 : _GEN_3844; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4877 = refillIDX_r & _GEN_12457 ? 1'h0 : _GEN_3845; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4878 = refillIDX_r & _GEN_12459 ? 1'h0 : _GEN_3846; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4879 = refillIDX_r & _GEN_12461 ? 1'h0 : _GEN_3847; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4880 = refillIDX_r & _GEN_12463 ? 1'h0 : _GEN_3848; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4881 = refillIDX_r & _GEN_12465 ? 1'h0 : _GEN_3849; // @[dcache.scala 424:{61,61}]
  wire  _GEN_4882 = refillIDX_r & _GEN_12467 ? 1'h0 : _GEN_3850; // @[dcache.scala 424:{61,61}]
  wire [20:0] _GEN_4883 = indexOnly ? _GEN_3851 : _GEN_4367; // @[dcache.scala 417:36]
  wire [20:0] _GEN_4884 = indexOnly ? _GEN_3852 : _GEN_4368; // @[dcache.scala 417:36]
  wire  _GEN_4885 = indexOnly ? _GEN_3853 : _GEN_4369; // @[dcache.scala 417:36]
  wire  _GEN_4886 = indexOnly ? _GEN_3854 : _GEN_4370; // @[dcache.scala 417:36]
  wire  _GEN_4887 = indexOnly ? _GEN_3855 : _GEN_4371; // @[dcache.scala 417:36]
  wire  _GEN_4888 = indexOnly ? _GEN_3856 : _GEN_4372; // @[dcache.scala 417:36]
  wire  _GEN_4889 = indexOnly ? _GEN_3857 : _GEN_4373; // @[dcache.scala 417:36]
  wire  _GEN_4890 = indexOnly ? _GEN_3858 : _GEN_4374; // @[dcache.scala 417:36]
  wire  _GEN_4891 = indexOnly ? _GEN_3859 : _GEN_4375; // @[dcache.scala 417:36]
  wire  _GEN_4892 = indexOnly ? _GEN_3860 : _GEN_4376; // @[dcache.scala 417:36]
  wire  _GEN_4893 = indexOnly ? _GEN_3861 : _GEN_4377; // @[dcache.scala 417:36]
  wire  _GEN_4894 = indexOnly ? _GEN_3862 : _GEN_4378; // @[dcache.scala 417:36]
  wire  _GEN_4895 = indexOnly ? _GEN_3863 : _GEN_4379; // @[dcache.scala 417:36]
  wire  _GEN_4896 = indexOnly ? _GEN_3864 : _GEN_4380; // @[dcache.scala 417:36]
  wire  _GEN_4897 = indexOnly ? _GEN_3865 : _GEN_4381; // @[dcache.scala 417:36]
  wire  _GEN_4898 = indexOnly ? _GEN_3866 : _GEN_4382; // @[dcache.scala 417:36]
  wire  _GEN_4899 = indexOnly ? _GEN_3867 : _GEN_4383; // @[dcache.scala 417:36]
  wire  _GEN_4900 = indexOnly ? _GEN_3868 : _GEN_4384; // @[dcache.scala 417:36]
  wire  _GEN_4901 = indexOnly ? _GEN_3869 : _GEN_4385; // @[dcache.scala 417:36]
  wire  _GEN_4902 = indexOnly ? _GEN_3870 : _GEN_4386; // @[dcache.scala 417:36]
  wire  _GEN_4903 = indexOnly ? _GEN_3871 : _GEN_4387; // @[dcache.scala 417:36]
  wire  _GEN_4904 = indexOnly ? _GEN_3872 : _GEN_4388; // @[dcache.scala 417:36]
  wire  _GEN_4905 = indexOnly ? _GEN_3873 : _GEN_4389; // @[dcache.scala 417:36]
  wire  _GEN_4906 = indexOnly ? _GEN_3874 : _GEN_4390; // @[dcache.scala 417:36]
  wire  _GEN_4907 = indexOnly ? _GEN_3875 : _GEN_4391; // @[dcache.scala 417:36]
  wire  _GEN_4908 = indexOnly ? _GEN_3876 : _GEN_4392; // @[dcache.scala 417:36]
  wire  _GEN_4909 = indexOnly ? _GEN_3877 : _GEN_4393; // @[dcache.scala 417:36]
  wire  _GEN_4910 = indexOnly ? _GEN_3878 : _GEN_4394; // @[dcache.scala 417:36]
  wire  _GEN_4911 = indexOnly ? _GEN_3879 : _GEN_4395; // @[dcache.scala 417:36]
  wire  _GEN_4912 = indexOnly ? _GEN_3880 : _GEN_4396; // @[dcache.scala 417:36]
  wire  _GEN_4913 = indexOnly ? _GEN_3881 : _GEN_4397; // @[dcache.scala 417:36]
  wire  _GEN_4914 = indexOnly ? _GEN_3882 : _GEN_4398; // @[dcache.scala 417:36]
  wire  _GEN_4915 = indexOnly ? _GEN_3883 : _GEN_4399; // @[dcache.scala 417:36]
  wire  _GEN_4916 = indexOnly ? _GEN_3884 : _GEN_4400; // @[dcache.scala 417:36]
  wire  _GEN_4917 = indexOnly ? _GEN_3885 : _GEN_4401; // @[dcache.scala 417:36]
  wire  _GEN_4918 = indexOnly ? _GEN_3886 : _GEN_4402; // @[dcache.scala 417:36]
  wire  _GEN_4919 = indexOnly ? _GEN_3887 : _GEN_4403; // @[dcache.scala 417:36]
  wire  _GEN_4920 = indexOnly ? _GEN_3888 : _GEN_4404; // @[dcache.scala 417:36]
  wire  _GEN_4921 = indexOnly ? _GEN_3889 : _GEN_4405; // @[dcache.scala 417:36]
  wire  _GEN_4922 = indexOnly ? _GEN_3890 : _GEN_4406; // @[dcache.scala 417:36]
  wire  _GEN_4923 = indexOnly ? _GEN_3891 : _GEN_4407; // @[dcache.scala 417:36]
  wire  _GEN_4924 = indexOnly ? _GEN_3892 : _GEN_4408; // @[dcache.scala 417:36]
  wire  _GEN_4925 = indexOnly ? _GEN_3893 : _GEN_4409; // @[dcache.scala 417:36]
  wire  _GEN_4926 = indexOnly ? _GEN_3894 : _GEN_4410; // @[dcache.scala 417:36]
  wire  _GEN_4927 = indexOnly ? _GEN_3895 : _GEN_4411; // @[dcache.scala 417:36]
  wire  _GEN_4928 = indexOnly ? _GEN_3896 : _GEN_4412; // @[dcache.scala 417:36]
  wire  _GEN_4929 = indexOnly ? _GEN_3897 : _GEN_4413; // @[dcache.scala 417:36]
  wire  _GEN_4930 = indexOnly ? _GEN_3898 : _GEN_4414; // @[dcache.scala 417:36]
  wire  _GEN_4931 = indexOnly ? _GEN_3899 : _GEN_4415; // @[dcache.scala 417:36]
  wire  _GEN_4932 = indexOnly ? _GEN_3900 : _GEN_4416; // @[dcache.scala 417:36]
  wire  _GEN_4933 = indexOnly ? _GEN_3901 : _GEN_4417; // @[dcache.scala 417:36]
  wire  _GEN_4934 = indexOnly ? _GEN_3902 : _GEN_4418; // @[dcache.scala 417:36]
  wire  _GEN_4935 = indexOnly ? _GEN_3903 : _GEN_4419; // @[dcache.scala 417:36]
  wire  _GEN_4936 = indexOnly ? _GEN_3904 : _GEN_4420; // @[dcache.scala 417:36]
  wire  _GEN_4937 = indexOnly ? _GEN_3905 : _GEN_4421; // @[dcache.scala 417:36]
  wire  _GEN_4938 = indexOnly ? _GEN_3906 : _GEN_4422; // @[dcache.scala 417:36]
  wire  _GEN_4939 = indexOnly ? _GEN_3907 : _GEN_4423; // @[dcache.scala 417:36]
  wire  _GEN_4940 = indexOnly ? _GEN_3908 : _GEN_4424; // @[dcache.scala 417:36]
  wire  _GEN_4941 = indexOnly ? _GEN_3909 : _GEN_4425; // @[dcache.scala 417:36]
  wire  _GEN_4942 = indexOnly ? _GEN_3910 : _GEN_4426; // @[dcache.scala 417:36]
  wire  _GEN_4943 = indexOnly ? _GEN_3911 : _GEN_4427; // @[dcache.scala 417:36]
  wire  _GEN_4944 = indexOnly ? _GEN_3912 : _GEN_4428; // @[dcache.scala 417:36]
  wire  _GEN_4945 = indexOnly ? _GEN_3913 : _GEN_4429; // @[dcache.scala 417:36]
  wire  _GEN_4946 = indexOnly ? _GEN_3914 : _GEN_4430; // @[dcache.scala 417:36]
  wire  _GEN_4947 = indexOnly ? _GEN_3915 : _GEN_4431; // @[dcache.scala 417:36]
  wire  _GEN_4948 = indexOnly ? _GEN_3916 : _GEN_4432; // @[dcache.scala 417:36]
  wire  _GEN_4949 = indexOnly ? _GEN_3917 : _GEN_4433; // @[dcache.scala 417:36]
  wire  _GEN_4950 = indexOnly ? _GEN_3918 : _GEN_4434; // @[dcache.scala 417:36]
  wire  _GEN_4951 = indexOnly ? _GEN_3919 : _GEN_4435; // @[dcache.scala 417:36]
  wire  _GEN_4952 = indexOnly ? _GEN_3920 : _GEN_4436; // @[dcache.scala 417:36]
  wire  _GEN_4953 = indexOnly ? _GEN_3921 : _GEN_4437; // @[dcache.scala 417:36]
  wire  _GEN_4954 = indexOnly ? _GEN_3922 : _GEN_4438; // @[dcache.scala 417:36]
  wire  _GEN_4955 = indexOnly ? _GEN_3923 : _GEN_4439; // @[dcache.scala 417:36]
  wire  _GEN_4956 = indexOnly ? _GEN_3924 : _GEN_4440; // @[dcache.scala 417:36]
  wire  _GEN_4957 = indexOnly ? _GEN_3925 : _GEN_4441; // @[dcache.scala 417:36]
  wire  _GEN_4958 = indexOnly ? _GEN_3926 : _GEN_4442; // @[dcache.scala 417:36]
  wire  _GEN_4959 = indexOnly ? _GEN_3927 : _GEN_4443; // @[dcache.scala 417:36]
  wire  _GEN_4960 = indexOnly ? _GEN_3928 : _GEN_4444; // @[dcache.scala 417:36]
  wire  _GEN_4961 = indexOnly ? _GEN_3929 : _GEN_4445; // @[dcache.scala 417:36]
  wire  _GEN_4962 = indexOnly ? _GEN_3930 : _GEN_4446; // @[dcache.scala 417:36]
  wire  _GEN_4963 = indexOnly ? _GEN_3931 : _GEN_4447; // @[dcache.scala 417:36]
  wire  _GEN_4964 = indexOnly ? _GEN_3932 : _GEN_4448; // @[dcache.scala 417:36]
  wire  _GEN_4965 = indexOnly ? _GEN_3933 : _GEN_4449; // @[dcache.scala 417:36]
  wire  _GEN_4966 = indexOnly ? _GEN_3934 : _GEN_4450; // @[dcache.scala 417:36]
  wire  _GEN_4967 = indexOnly ? _GEN_3935 : _GEN_4451; // @[dcache.scala 417:36]
  wire  _GEN_4968 = indexOnly ? _GEN_3936 : _GEN_4452; // @[dcache.scala 417:36]
  wire  _GEN_4969 = indexOnly ? _GEN_3937 : _GEN_4453; // @[dcache.scala 417:36]
  wire  _GEN_4970 = indexOnly ? _GEN_3938 : _GEN_4454; // @[dcache.scala 417:36]
  wire  _GEN_4971 = indexOnly ? _GEN_3939 : _GEN_4455; // @[dcache.scala 417:36]
  wire  _GEN_4972 = indexOnly ? _GEN_3940 : _GEN_4456; // @[dcache.scala 417:36]
  wire  _GEN_4973 = indexOnly ? _GEN_3941 : _GEN_4457; // @[dcache.scala 417:36]
  wire  _GEN_4974 = indexOnly ? _GEN_3942 : _GEN_4458; // @[dcache.scala 417:36]
  wire  _GEN_4975 = indexOnly ? _GEN_3943 : _GEN_4459; // @[dcache.scala 417:36]
  wire  _GEN_4976 = indexOnly ? _GEN_3944 : _GEN_4460; // @[dcache.scala 417:36]
  wire  _GEN_4977 = indexOnly ? _GEN_3945 : _GEN_4461; // @[dcache.scala 417:36]
  wire  _GEN_4978 = indexOnly ? _GEN_3946 : _GEN_4462; // @[dcache.scala 417:36]
  wire  _GEN_4979 = indexOnly ? _GEN_3947 : _GEN_4463; // @[dcache.scala 417:36]
  wire  _GEN_4980 = indexOnly ? _GEN_3948 : _GEN_4464; // @[dcache.scala 417:36]
  wire  _GEN_4981 = indexOnly ? _GEN_3949 : _GEN_4465; // @[dcache.scala 417:36]
  wire  _GEN_4982 = indexOnly ? _GEN_3950 : _GEN_4466; // @[dcache.scala 417:36]
  wire  _GEN_4983 = indexOnly ? _GEN_3951 : _GEN_4467; // @[dcache.scala 417:36]
  wire  _GEN_4984 = indexOnly ? _GEN_3952 : _GEN_4468; // @[dcache.scala 417:36]
  wire  _GEN_4985 = indexOnly ? _GEN_3953 : _GEN_4469; // @[dcache.scala 417:36]
  wire  _GEN_4986 = indexOnly ? _GEN_3954 : _GEN_4470; // @[dcache.scala 417:36]
  wire  _GEN_4987 = indexOnly ? _GEN_3955 : _GEN_4471; // @[dcache.scala 417:36]
  wire  _GEN_4988 = indexOnly ? _GEN_3956 : _GEN_4472; // @[dcache.scala 417:36]
  wire  _GEN_4989 = indexOnly ? _GEN_3957 : _GEN_4473; // @[dcache.scala 417:36]
  wire  _GEN_4990 = indexOnly ? _GEN_3958 : _GEN_4474; // @[dcache.scala 417:36]
  wire  _GEN_4991 = indexOnly ? _GEN_3959 : _GEN_4475; // @[dcache.scala 417:36]
  wire  _GEN_4992 = indexOnly ? _GEN_3960 : _GEN_4476; // @[dcache.scala 417:36]
  wire  _GEN_4993 = indexOnly ? _GEN_3961 : _GEN_4477; // @[dcache.scala 417:36]
  wire  _GEN_4994 = indexOnly ? _GEN_3962 : _GEN_4478; // @[dcache.scala 417:36]
  wire  _GEN_4995 = indexOnly ? _GEN_3963 : _GEN_4479; // @[dcache.scala 417:36]
  wire  _GEN_4996 = indexOnly ? _GEN_3964 : _GEN_4480; // @[dcache.scala 417:36]
  wire  _GEN_4997 = indexOnly ? _GEN_3965 : _GEN_4481; // @[dcache.scala 417:36]
  wire  _GEN_4998 = indexOnly ? _GEN_3966 : _GEN_4482; // @[dcache.scala 417:36]
  wire  _GEN_4999 = indexOnly ? _GEN_3967 : _GEN_4483; // @[dcache.scala 417:36]
  wire  _GEN_5000 = indexOnly ? _GEN_3968 : _GEN_4484; // @[dcache.scala 417:36]
  wire  _GEN_5001 = indexOnly ? _GEN_3969 : _GEN_4485; // @[dcache.scala 417:36]
  wire  _GEN_5002 = indexOnly ? _GEN_3970 : _GEN_4486; // @[dcache.scala 417:36]
  wire  _GEN_5003 = indexOnly ? _GEN_3971 : _GEN_4487; // @[dcache.scala 417:36]
  wire  _GEN_5004 = indexOnly ? _GEN_3972 : _GEN_4488; // @[dcache.scala 417:36]
  wire  _GEN_5005 = indexOnly ? _GEN_3973 : _GEN_4489; // @[dcache.scala 417:36]
  wire  _GEN_5006 = indexOnly ? _GEN_3974 : _GEN_4490; // @[dcache.scala 417:36]
  wire  _GEN_5007 = indexOnly ? _GEN_3975 : _GEN_4491; // @[dcache.scala 417:36]
  wire  _GEN_5008 = indexOnly ? _GEN_3976 : _GEN_4492; // @[dcache.scala 417:36]
  wire  _GEN_5009 = indexOnly ? _GEN_3977 : _GEN_4493; // @[dcache.scala 417:36]
  wire  _GEN_5010 = indexOnly ? _GEN_3978 : _GEN_4494; // @[dcache.scala 417:36]
  wire  _GEN_5011 = indexOnly ? _GEN_3979 : _GEN_4495; // @[dcache.scala 417:36]
  wire  _GEN_5012 = indexOnly ? _GEN_3980 : _GEN_4496; // @[dcache.scala 417:36]
  wire  _GEN_5013 = indexOnly ? _GEN_3981 : _GEN_4497; // @[dcache.scala 417:36]
  wire  _GEN_5014 = indexOnly ? _GEN_3982 : _GEN_4498; // @[dcache.scala 417:36]
  wire  _GEN_5015 = indexOnly ? _GEN_3983 : _GEN_4499; // @[dcache.scala 417:36]
  wire  _GEN_5016 = indexOnly ? _GEN_3984 : _GEN_4500; // @[dcache.scala 417:36]
  wire  _GEN_5017 = indexOnly ? _GEN_3985 : _GEN_4501; // @[dcache.scala 417:36]
  wire  _GEN_5018 = indexOnly ? _GEN_3986 : _GEN_4502; // @[dcache.scala 417:36]
  wire  _GEN_5019 = indexOnly ? _GEN_3987 : _GEN_4503; // @[dcache.scala 417:36]
  wire  _GEN_5020 = indexOnly ? _GEN_3988 : _GEN_4504; // @[dcache.scala 417:36]
  wire  _GEN_5021 = indexOnly ? _GEN_3989 : _GEN_4505; // @[dcache.scala 417:36]
  wire  _GEN_5022 = indexOnly ? _GEN_3990 : _GEN_4506; // @[dcache.scala 417:36]
  wire  _GEN_5023 = indexOnly ? _GEN_3991 : _GEN_4507; // @[dcache.scala 417:36]
  wire  _GEN_5024 = indexOnly ? _GEN_3992 : _GEN_4508; // @[dcache.scala 417:36]
  wire  _GEN_5025 = indexOnly ? _GEN_3993 : _GEN_4509; // @[dcache.scala 417:36]
  wire  _GEN_5026 = indexOnly ? _GEN_3994 : _GEN_4510; // @[dcache.scala 417:36]
  wire  _GEN_5027 = indexOnly ? _GEN_3995 : _GEN_4511; // @[dcache.scala 417:36]
  wire  _GEN_5028 = indexOnly ? _GEN_3996 : _GEN_4512; // @[dcache.scala 417:36]
  wire  _GEN_5029 = indexOnly ? _GEN_3997 : _GEN_4513; // @[dcache.scala 417:36]
  wire  _GEN_5030 = indexOnly ? _GEN_3998 : _GEN_4514; // @[dcache.scala 417:36]
  wire  _GEN_5031 = indexOnly ? _GEN_3999 : _GEN_4515; // @[dcache.scala 417:36]
  wire  _GEN_5032 = indexOnly ? _GEN_4000 : _GEN_4516; // @[dcache.scala 417:36]
  wire  _GEN_5033 = indexOnly ? _GEN_4001 : _GEN_4517; // @[dcache.scala 417:36]
  wire  _GEN_5034 = indexOnly ? _GEN_4002 : _GEN_4518; // @[dcache.scala 417:36]
  wire  _GEN_5035 = indexOnly ? _GEN_4003 : _GEN_4519; // @[dcache.scala 417:36]
  wire  _GEN_5036 = indexOnly ? _GEN_4004 : _GEN_4520; // @[dcache.scala 417:36]
  wire  _GEN_5037 = indexOnly ? _GEN_4005 : _GEN_4521; // @[dcache.scala 417:36]
  wire  _GEN_5038 = indexOnly ? _GEN_4006 : _GEN_4522; // @[dcache.scala 417:36]
  wire  _GEN_5039 = indexOnly ? _GEN_4007 : _GEN_4523; // @[dcache.scala 417:36]
  wire  _GEN_5040 = indexOnly ? _GEN_4008 : _GEN_4524; // @[dcache.scala 417:36]
  wire  _GEN_5041 = indexOnly ? _GEN_4009 : _GEN_4525; // @[dcache.scala 417:36]
  wire  _GEN_5042 = indexOnly ? _GEN_4010 : _GEN_4526; // @[dcache.scala 417:36]
  wire  _GEN_5043 = indexOnly ? _GEN_4011 : _GEN_4527; // @[dcache.scala 417:36]
  wire  _GEN_5044 = indexOnly ? _GEN_4012 : _GEN_4528; // @[dcache.scala 417:36]
  wire  _GEN_5045 = indexOnly ? _GEN_4013 : _GEN_4529; // @[dcache.scala 417:36]
  wire  _GEN_5046 = indexOnly ? _GEN_4014 : _GEN_4530; // @[dcache.scala 417:36]
  wire  _GEN_5047 = indexOnly ? _GEN_4015 : _GEN_4531; // @[dcache.scala 417:36]
  wire  _GEN_5048 = indexOnly ? _GEN_4016 : _GEN_4532; // @[dcache.scala 417:36]
  wire  _GEN_5049 = indexOnly ? _GEN_4017 : _GEN_4533; // @[dcache.scala 417:36]
  wire  _GEN_5050 = indexOnly ? _GEN_4018 : _GEN_4534; // @[dcache.scala 417:36]
  wire  _GEN_5051 = indexOnly ? _GEN_4019 : _GEN_4535; // @[dcache.scala 417:36]
  wire  _GEN_5052 = indexOnly ? _GEN_4020 : _GEN_4536; // @[dcache.scala 417:36]
  wire  _GEN_5053 = indexOnly ? _GEN_4021 : _GEN_4537; // @[dcache.scala 417:36]
  wire  _GEN_5054 = indexOnly ? _GEN_4022 : _GEN_4538; // @[dcache.scala 417:36]
  wire  _GEN_5055 = indexOnly ? _GEN_4023 : _GEN_4539; // @[dcache.scala 417:36]
  wire  _GEN_5056 = indexOnly ? _GEN_4024 : _GEN_4540; // @[dcache.scala 417:36]
  wire  _GEN_5057 = indexOnly ? _GEN_4025 : _GEN_4541; // @[dcache.scala 417:36]
  wire  _GEN_5058 = indexOnly ? _GEN_4026 : _GEN_4542; // @[dcache.scala 417:36]
  wire  _GEN_5059 = indexOnly ? _GEN_4027 : _GEN_4543; // @[dcache.scala 417:36]
  wire  _GEN_5060 = indexOnly ? _GEN_4028 : _GEN_4544; // @[dcache.scala 417:36]
  wire  _GEN_5061 = indexOnly ? _GEN_4029 : _GEN_4545; // @[dcache.scala 417:36]
  wire  _GEN_5062 = indexOnly ? _GEN_4030 : _GEN_4546; // @[dcache.scala 417:36]
  wire  _GEN_5063 = indexOnly ? _GEN_4031 : _GEN_4547; // @[dcache.scala 417:36]
  wire  _GEN_5064 = indexOnly ? _GEN_4032 : _GEN_4548; // @[dcache.scala 417:36]
  wire  _GEN_5065 = indexOnly ? _GEN_4033 : _GEN_4549; // @[dcache.scala 417:36]
  wire  _GEN_5066 = indexOnly ? _GEN_4034 : _GEN_4550; // @[dcache.scala 417:36]
  wire  _GEN_5067 = indexOnly ? _GEN_4035 : _GEN_4551; // @[dcache.scala 417:36]
  wire  _GEN_5068 = indexOnly ? _GEN_4036 : _GEN_4552; // @[dcache.scala 417:36]
  wire  _GEN_5069 = indexOnly ? _GEN_4037 : _GEN_4553; // @[dcache.scala 417:36]
  wire  _GEN_5070 = indexOnly ? _GEN_4038 : _GEN_4554; // @[dcache.scala 417:36]
  wire  _GEN_5071 = indexOnly ? _GEN_4039 : _GEN_4555; // @[dcache.scala 417:36]
  wire  _GEN_5072 = indexOnly ? _GEN_4040 : _GEN_4556; // @[dcache.scala 417:36]
  wire  _GEN_5073 = indexOnly ? _GEN_4041 : _GEN_4557; // @[dcache.scala 417:36]
  wire  _GEN_5074 = indexOnly ? _GEN_4042 : _GEN_4558; // @[dcache.scala 417:36]
  wire  _GEN_5075 = indexOnly ? _GEN_4043 : _GEN_4559; // @[dcache.scala 417:36]
  wire  _GEN_5076 = indexOnly ? _GEN_4044 : _GEN_4560; // @[dcache.scala 417:36]
  wire  _GEN_5077 = indexOnly ? _GEN_4045 : _GEN_4561; // @[dcache.scala 417:36]
  wire  _GEN_5078 = indexOnly ? _GEN_4046 : _GEN_4562; // @[dcache.scala 417:36]
  wire  _GEN_5079 = indexOnly ? _GEN_4047 : _GEN_4563; // @[dcache.scala 417:36]
  wire  _GEN_5080 = indexOnly ? _GEN_4048 : _GEN_4564; // @[dcache.scala 417:36]
  wire  _GEN_5081 = indexOnly ? _GEN_4049 : _GEN_4565; // @[dcache.scala 417:36]
  wire  _GEN_5082 = indexOnly ? _GEN_4050 : _GEN_4566; // @[dcache.scala 417:36]
  wire  _GEN_5083 = indexOnly ? _GEN_4051 : _GEN_4567; // @[dcache.scala 417:36]
  wire  _GEN_5084 = indexOnly ? _GEN_4052 : _GEN_4568; // @[dcache.scala 417:36]
  wire  _GEN_5085 = indexOnly ? _GEN_4053 : _GEN_4569; // @[dcache.scala 417:36]
  wire  _GEN_5086 = indexOnly ? _GEN_4054 : _GEN_4570; // @[dcache.scala 417:36]
  wire  _GEN_5087 = indexOnly ? _GEN_4055 : _GEN_4571; // @[dcache.scala 417:36]
  wire  _GEN_5088 = indexOnly ? _GEN_4056 : _GEN_4572; // @[dcache.scala 417:36]
  wire  _GEN_5089 = indexOnly ? _GEN_4057 : _GEN_4573; // @[dcache.scala 417:36]
  wire  _GEN_5090 = indexOnly ? _GEN_4058 : _GEN_4574; // @[dcache.scala 417:36]
  wire  _GEN_5091 = indexOnly ? _GEN_4059 : _GEN_4575; // @[dcache.scala 417:36]
  wire  _GEN_5092 = indexOnly ? _GEN_4060 : _GEN_4576; // @[dcache.scala 417:36]
  wire  _GEN_5093 = indexOnly ? _GEN_4061 : _GEN_4577; // @[dcache.scala 417:36]
  wire  _GEN_5094 = indexOnly ? _GEN_4062 : _GEN_4578; // @[dcache.scala 417:36]
  wire  _GEN_5095 = indexOnly ? _GEN_4063 : _GEN_4579; // @[dcache.scala 417:36]
  wire  _GEN_5096 = indexOnly ? _GEN_4064 : _GEN_4580; // @[dcache.scala 417:36]
  wire  _GEN_5097 = indexOnly ? _GEN_4065 : _GEN_4581; // @[dcache.scala 417:36]
  wire  _GEN_5098 = indexOnly ? _GEN_4066 : _GEN_4582; // @[dcache.scala 417:36]
  wire  _GEN_5099 = indexOnly ? _GEN_4067 : _GEN_4583; // @[dcache.scala 417:36]
  wire  _GEN_5100 = indexOnly ? _GEN_4068 : _GEN_4584; // @[dcache.scala 417:36]
  wire  _GEN_5101 = indexOnly ? _GEN_4069 : _GEN_4585; // @[dcache.scala 417:36]
  wire  _GEN_5102 = indexOnly ? _GEN_4070 : _GEN_4586; // @[dcache.scala 417:36]
  wire  _GEN_5103 = indexOnly ? _GEN_4071 : _GEN_4587; // @[dcache.scala 417:36]
  wire  _GEN_5104 = indexOnly ? _GEN_4072 : _GEN_4588; // @[dcache.scala 417:36]
  wire  _GEN_5105 = indexOnly ? _GEN_4073 : _GEN_4589; // @[dcache.scala 417:36]
  wire  _GEN_5106 = indexOnly ? _GEN_4074 : _GEN_4590; // @[dcache.scala 417:36]
  wire  _GEN_5107 = indexOnly ? _GEN_4075 : _GEN_4591; // @[dcache.scala 417:36]
  wire  _GEN_5108 = indexOnly ? _GEN_4076 : _GEN_4592; // @[dcache.scala 417:36]
  wire  _GEN_5109 = indexOnly ? _GEN_4077 : _GEN_4593; // @[dcache.scala 417:36]
  wire  _GEN_5110 = indexOnly ? _GEN_4078 : _GEN_4594; // @[dcache.scala 417:36]
  wire  _GEN_5111 = indexOnly ? _GEN_4079 : _GEN_4595; // @[dcache.scala 417:36]
  wire  _GEN_5112 = indexOnly ? _GEN_4080 : _GEN_4596; // @[dcache.scala 417:36]
  wire  _GEN_5113 = indexOnly ? _GEN_4081 : _GEN_4597; // @[dcache.scala 417:36]
  wire  _GEN_5114 = indexOnly ? _GEN_4082 : _GEN_4598; // @[dcache.scala 417:36]
  wire  _GEN_5115 = indexOnly ? _GEN_4083 : _GEN_4599; // @[dcache.scala 417:36]
  wire  _GEN_5116 = indexOnly ? _GEN_4084 : _GEN_4600; // @[dcache.scala 417:36]
  wire  _GEN_5117 = indexOnly ? _GEN_4085 : _GEN_4601; // @[dcache.scala 417:36]
  wire  _GEN_5118 = indexOnly ? _GEN_4086 : _GEN_4602; // @[dcache.scala 417:36]
  wire  _GEN_5119 = indexOnly ? _GEN_4087 : _GEN_4603; // @[dcache.scala 417:36]
  wire  _GEN_5120 = indexOnly ? _GEN_4088 : _GEN_4604; // @[dcache.scala 417:36]
  wire  _GEN_5121 = indexOnly ? _GEN_4089 : _GEN_4605; // @[dcache.scala 417:36]
  wire  _GEN_5122 = indexOnly ? _GEN_4090 : _GEN_4606; // @[dcache.scala 417:36]
  wire  _GEN_5123 = indexOnly ? _GEN_4091 : _GEN_4607; // @[dcache.scala 417:36]
  wire  _GEN_5124 = indexOnly ? _GEN_4092 : _GEN_4608; // @[dcache.scala 417:36]
  wire  _GEN_5125 = indexOnly ? _GEN_4093 : _GEN_4609; // @[dcache.scala 417:36]
  wire  _GEN_5126 = indexOnly ? _GEN_4094 : _GEN_4610; // @[dcache.scala 417:36]
  wire  _GEN_5127 = indexOnly ? _GEN_4095 : _GEN_4611; // @[dcache.scala 417:36]
  wire  _GEN_5128 = indexOnly ? _GEN_4096 : _GEN_4612; // @[dcache.scala 417:36]
  wire  _GEN_5129 = indexOnly ? _GEN_4097 : _GEN_4613; // @[dcache.scala 417:36]
  wire  _GEN_5130 = indexOnly ? _GEN_4098 : _GEN_4614; // @[dcache.scala 417:36]
  wire  _GEN_5131 = indexOnly ? _GEN_4099 : _GEN_4615; // @[dcache.scala 417:36]
  wire  _GEN_5132 = indexOnly ? _GEN_4100 : _GEN_4616; // @[dcache.scala 417:36]
  wire  _GEN_5133 = indexOnly ? _GEN_4101 : _GEN_4617; // @[dcache.scala 417:36]
  wire  _GEN_5134 = indexOnly ? _GEN_4102 : _GEN_4618; // @[dcache.scala 417:36]
  wire  _GEN_5135 = indexOnly ? _GEN_4103 : _GEN_4619; // @[dcache.scala 417:36]
  wire  _GEN_5136 = indexOnly ? _GEN_4104 : _GEN_4620; // @[dcache.scala 417:36]
  wire  _GEN_5137 = indexOnly ? _GEN_4105 : _GEN_4621; // @[dcache.scala 417:36]
  wire  _GEN_5138 = indexOnly ? _GEN_4106 : _GEN_4622; // @[dcache.scala 417:36]
  wire  _GEN_5139 = indexOnly ? _GEN_4107 : _GEN_4623; // @[dcache.scala 417:36]
  wire  _GEN_5140 = indexOnly ? _GEN_4108 : _GEN_4624; // @[dcache.scala 417:36]
  wire  _GEN_5141 = indexOnly ? _GEN_4109 : _GEN_4625; // @[dcache.scala 417:36]
  wire  _GEN_5142 = indexOnly ? _GEN_4110 : _GEN_4626; // @[dcache.scala 417:36]
  wire  _GEN_5143 = indexOnly ? _GEN_4111 : _GEN_4627; // @[dcache.scala 417:36]
  wire  _GEN_5144 = indexOnly ? _GEN_4112 : _GEN_4628; // @[dcache.scala 417:36]
  wire  _GEN_5145 = indexOnly ? _GEN_4113 : _GEN_4629; // @[dcache.scala 417:36]
  wire  _GEN_5146 = indexOnly ? _GEN_4114 : _GEN_4630; // @[dcache.scala 417:36]
  wire  _GEN_5147 = indexOnly ? _GEN_4115 : _GEN_4631; // @[dcache.scala 417:36]
  wire  _GEN_5148 = indexOnly ? _GEN_4116 : _GEN_4632; // @[dcache.scala 417:36]
  wire  _GEN_5149 = indexOnly ? _GEN_4117 : _GEN_4633; // @[dcache.scala 417:36]
  wire  _GEN_5150 = indexOnly ? _GEN_4118 : _GEN_4634; // @[dcache.scala 417:36]
  wire  _GEN_5151 = indexOnly ? _GEN_4119 : _GEN_4635; // @[dcache.scala 417:36]
  wire  _GEN_5152 = indexOnly ? _GEN_4120 : _GEN_4636; // @[dcache.scala 417:36]
  wire  _GEN_5153 = indexOnly ? _GEN_4121 : _GEN_4637; // @[dcache.scala 417:36]
  wire  _GEN_5154 = indexOnly ? _GEN_4122 : _GEN_4638; // @[dcache.scala 417:36]
  wire  _GEN_5155 = indexOnly ? _GEN_4123 : _GEN_4639; // @[dcache.scala 417:36]
  wire  _GEN_5156 = indexOnly ? _GEN_4124 : _GEN_4640; // @[dcache.scala 417:36]
  wire  _GEN_5157 = indexOnly ? _GEN_4125 : _GEN_4641; // @[dcache.scala 417:36]
  wire  _GEN_5158 = indexOnly ? _GEN_4126 : _GEN_4642; // @[dcache.scala 417:36]
  wire  _GEN_5159 = indexOnly ? _GEN_4127 : _GEN_4643; // @[dcache.scala 417:36]
  wire  _GEN_5160 = indexOnly ? _GEN_4128 : _GEN_4644; // @[dcache.scala 417:36]
  wire  _GEN_5161 = indexOnly ? _GEN_4129 : _GEN_4645; // @[dcache.scala 417:36]
  wire  _GEN_5162 = indexOnly ? _GEN_4130 : _GEN_4646; // @[dcache.scala 417:36]
  wire  _GEN_5163 = indexOnly ? _GEN_4131 : _GEN_4647; // @[dcache.scala 417:36]
  wire  _GEN_5164 = indexOnly ? _GEN_4132 : _GEN_4648; // @[dcache.scala 417:36]
  wire  _GEN_5165 = indexOnly ? _GEN_4133 : _GEN_4649; // @[dcache.scala 417:36]
  wire  _GEN_5166 = indexOnly ? _GEN_4134 : _GEN_4650; // @[dcache.scala 417:36]
  wire  _GEN_5167 = indexOnly ? _GEN_4135 : _GEN_4651; // @[dcache.scala 417:36]
  wire  _GEN_5168 = indexOnly ? _GEN_4136 : _GEN_4652; // @[dcache.scala 417:36]
  wire  _GEN_5169 = indexOnly ? _GEN_4137 : _GEN_4653; // @[dcache.scala 417:36]
  wire  _GEN_5170 = indexOnly ? _GEN_4138 : _GEN_4654; // @[dcache.scala 417:36]
  wire  _GEN_5171 = indexOnly ? _GEN_4139 : _GEN_4655; // @[dcache.scala 417:36]
  wire  _GEN_5172 = indexOnly ? _GEN_4140 : _GEN_4656; // @[dcache.scala 417:36]
  wire  _GEN_5173 = indexOnly ? _GEN_4141 : _GEN_4657; // @[dcache.scala 417:36]
  wire  _GEN_5174 = indexOnly ? _GEN_4142 : _GEN_4658; // @[dcache.scala 417:36]
  wire  _GEN_5175 = indexOnly ? _GEN_4143 : _GEN_4659; // @[dcache.scala 417:36]
  wire  _GEN_5176 = indexOnly ? _GEN_4144 : _GEN_4660; // @[dcache.scala 417:36]
  wire  _GEN_5177 = indexOnly ? _GEN_4145 : _GEN_4661; // @[dcache.scala 417:36]
  wire  _GEN_5178 = indexOnly ? _GEN_4146 : _GEN_4662; // @[dcache.scala 417:36]
  wire  _GEN_5179 = indexOnly ? _GEN_4147 : _GEN_4663; // @[dcache.scala 417:36]
  wire  _GEN_5180 = indexOnly ? _GEN_4148 : _GEN_4664; // @[dcache.scala 417:36]
  wire  _GEN_5181 = indexOnly ? _GEN_4149 : _GEN_4665; // @[dcache.scala 417:36]
  wire  _GEN_5182 = indexOnly ? _GEN_4150 : _GEN_4666; // @[dcache.scala 417:36]
  wire  _GEN_5183 = indexOnly ? _GEN_4151 : _GEN_4667; // @[dcache.scala 417:36]
  wire  _GEN_5184 = indexOnly ? _GEN_4152 : _GEN_4668; // @[dcache.scala 417:36]
  wire  _GEN_5185 = indexOnly ? _GEN_4153 : _GEN_4669; // @[dcache.scala 417:36]
  wire  _GEN_5186 = indexOnly ? _GEN_4154 : _GEN_4670; // @[dcache.scala 417:36]
  wire  _GEN_5187 = indexOnly ? _GEN_4155 : _GEN_4671; // @[dcache.scala 417:36]
  wire  _GEN_5188 = indexOnly ? _GEN_4156 : _GEN_4672; // @[dcache.scala 417:36]
  wire  _GEN_5189 = indexOnly ? _GEN_4157 : _GEN_4673; // @[dcache.scala 417:36]
  wire  _GEN_5190 = indexOnly ? _GEN_4158 : _GEN_4674; // @[dcache.scala 417:36]
  wire  _GEN_5191 = indexOnly ? _GEN_4159 : _GEN_4675; // @[dcache.scala 417:36]
  wire  _GEN_5192 = indexOnly ? _GEN_4160 : _GEN_4676; // @[dcache.scala 417:36]
  wire  _GEN_5193 = indexOnly ? _GEN_4161 : _GEN_4677; // @[dcache.scala 417:36]
  wire  _GEN_5194 = indexOnly ? _GEN_4162 : _GEN_4678; // @[dcache.scala 417:36]
  wire  _GEN_5195 = indexOnly ? _GEN_4163 : _GEN_4679; // @[dcache.scala 417:36]
  wire  _GEN_5196 = indexOnly ? _GEN_4164 : _GEN_4680; // @[dcache.scala 417:36]
  wire  _GEN_5197 = indexOnly ? _GEN_4165 : _GEN_4681; // @[dcache.scala 417:36]
  wire  _GEN_5198 = indexOnly ? _GEN_4166 : _GEN_4682; // @[dcache.scala 417:36]
  wire  _GEN_5199 = indexOnly ? _GEN_4167 : _GEN_4683; // @[dcache.scala 417:36]
  wire  _GEN_5200 = indexOnly ? _GEN_4168 : _GEN_4684; // @[dcache.scala 417:36]
  wire  _GEN_5201 = indexOnly ? _GEN_4169 : _GEN_4685; // @[dcache.scala 417:36]
  wire  _GEN_5202 = indexOnly ? _GEN_4170 : _GEN_4686; // @[dcache.scala 417:36]
  wire  _GEN_5203 = indexOnly ? _GEN_4171 : _GEN_4687; // @[dcache.scala 417:36]
  wire  _GEN_5204 = indexOnly ? _GEN_4172 : _GEN_4688; // @[dcache.scala 417:36]
  wire  _GEN_5205 = indexOnly ? _GEN_4173 : _GEN_4689; // @[dcache.scala 417:36]
  wire  _GEN_5206 = indexOnly ? _GEN_4174 : _GEN_4690; // @[dcache.scala 417:36]
  wire  _GEN_5207 = indexOnly ? _GEN_4175 : _GEN_4691; // @[dcache.scala 417:36]
  wire  _GEN_5208 = indexOnly ? _GEN_4176 : _GEN_4692; // @[dcache.scala 417:36]
  wire  _GEN_5209 = indexOnly ? _GEN_4177 : _GEN_4693; // @[dcache.scala 417:36]
  wire  _GEN_5210 = indexOnly ? _GEN_4178 : _GEN_4694; // @[dcache.scala 417:36]
  wire  _GEN_5211 = indexOnly ? _GEN_4179 : _GEN_4695; // @[dcache.scala 417:36]
  wire  _GEN_5212 = indexOnly ? _GEN_4180 : _GEN_4696; // @[dcache.scala 417:36]
  wire  _GEN_5213 = indexOnly ? _GEN_4181 : _GEN_4697; // @[dcache.scala 417:36]
  wire  _GEN_5214 = indexOnly ? _GEN_4182 : _GEN_4698; // @[dcache.scala 417:36]
  wire  _GEN_5215 = indexOnly ? _GEN_4183 : _GEN_4699; // @[dcache.scala 417:36]
  wire  _GEN_5216 = indexOnly ? _GEN_4184 : _GEN_4700; // @[dcache.scala 417:36]
  wire  _GEN_5217 = indexOnly ? _GEN_4185 : _GEN_4701; // @[dcache.scala 417:36]
  wire  _GEN_5218 = indexOnly ? _GEN_4186 : _GEN_4702; // @[dcache.scala 417:36]
  wire  _GEN_5219 = indexOnly ? _GEN_4187 : _GEN_4703; // @[dcache.scala 417:36]
  wire  _GEN_5220 = indexOnly ? _GEN_4188 : _GEN_4704; // @[dcache.scala 417:36]
  wire  _GEN_5221 = indexOnly ? _GEN_4189 : _GEN_4705; // @[dcache.scala 417:36]
  wire  _GEN_5222 = indexOnly ? _GEN_4190 : _GEN_4706; // @[dcache.scala 417:36]
  wire  _GEN_5223 = indexOnly ? _GEN_4191 : _GEN_4707; // @[dcache.scala 417:36]
  wire  _GEN_5224 = indexOnly ? _GEN_4192 : _GEN_4708; // @[dcache.scala 417:36]
  wire  _GEN_5225 = indexOnly ? _GEN_4193 : _GEN_4709; // @[dcache.scala 417:36]
  wire  _GEN_5226 = indexOnly ? _GEN_4194 : _GEN_4710; // @[dcache.scala 417:36]
  wire  _GEN_5227 = indexOnly ? _GEN_4195 : _GEN_4711; // @[dcache.scala 417:36]
  wire  _GEN_5228 = indexOnly ? _GEN_4196 : _GEN_4712; // @[dcache.scala 417:36]
  wire  _GEN_5229 = indexOnly ? _GEN_4197 : _GEN_4713; // @[dcache.scala 417:36]
  wire  _GEN_5230 = indexOnly ? _GEN_4198 : _GEN_4714; // @[dcache.scala 417:36]
  wire  _GEN_5231 = indexOnly ? _GEN_4199 : _GEN_4715; // @[dcache.scala 417:36]
  wire  _GEN_5232 = indexOnly ? _GEN_4200 : _GEN_4716; // @[dcache.scala 417:36]
  wire  _GEN_5233 = indexOnly ? _GEN_4201 : _GEN_4717; // @[dcache.scala 417:36]
  wire  _GEN_5234 = indexOnly ? _GEN_4202 : _GEN_4718; // @[dcache.scala 417:36]
  wire  _GEN_5235 = indexOnly ? _GEN_4203 : _GEN_4719; // @[dcache.scala 417:36]
  wire  _GEN_5236 = indexOnly ? _GEN_4204 : _GEN_4720; // @[dcache.scala 417:36]
  wire  _GEN_5237 = indexOnly ? _GEN_4205 : _GEN_4721; // @[dcache.scala 417:36]
  wire  _GEN_5238 = indexOnly ? _GEN_4206 : _GEN_4722; // @[dcache.scala 417:36]
  wire  _GEN_5239 = indexOnly ? _GEN_4207 : _GEN_4723; // @[dcache.scala 417:36]
  wire  _GEN_5240 = indexOnly ? _GEN_4208 : _GEN_4724; // @[dcache.scala 417:36]
  wire  _GEN_5241 = indexOnly ? _GEN_4209 : _GEN_4725; // @[dcache.scala 417:36]
  wire  _GEN_5242 = indexOnly ? _GEN_4210 : _GEN_4726; // @[dcache.scala 417:36]
  wire  _GEN_5243 = indexOnly ? _GEN_4211 : _GEN_4727; // @[dcache.scala 417:36]
  wire  _GEN_5244 = indexOnly ? _GEN_4212 : _GEN_4728; // @[dcache.scala 417:36]
  wire  _GEN_5245 = indexOnly ? _GEN_4213 : _GEN_4729; // @[dcache.scala 417:36]
  wire  _GEN_5246 = indexOnly ? _GEN_4214 : _GEN_4730; // @[dcache.scala 417:36]
  wire  _GEN_5247 = indexOnly ? _GEN_4215 : _GEN_4731; // @[dcache.scala 417:36]
  wire  _GEN_5248 = indexOnly ? _GEN_4216 : _GEN_4732; // @[dcache.scala 417:36]
  wire  _GEN_5249 = indexOnly ? _GEN_4217 : _GEN_4733; // @[dcache.scala 417:36]
  wire  _GEN_5250 = indexOnly ? _GEN_4218 : _GEN_4734; // @[dcache.scala 417:36]
  wire  _GEN_5251 = indexOnly ? _GEN_4219 : _GEN_4735; // @[dcache.scala 417:36]
  wire  _GEN_5252 = indexOnly ? _GEN_4220 : _GEN_4736; // @[dcache.scala 417:36]
  wire  _GEN_5253 = indexOnly ? _GEN_4221 : _GEN_4737; // @[dcache.scala 417:36]
  wire  _GEN_5254 = indexOnly ? _GEN_4222 : _GEN_4738; // @[dcache.scala 417:36]
  wire  _GEN_5255 = indexOnly ? _GEN_4223 : _GEN_4739; // @[dcache.scala 417:36]
  wire  _GEN_5256 = indexOnly ? _GEN_4224 : _GEN_4740; // @[dcache.scala 417:36]
  wire  _GEN_5257 = indexOnly ? _GEN_4225 : _GEN_4741; // @[dcache.scala 417:36]
  wire  _GEN_5258 = indexOnly ? _GEN_4226 : _GEN_4742; // @[dcache.scala 417:36]
  wire  _GEN_5259 = indexOnly ? _GEN_4227 : _GEN_4743; // @[dcache.scala 417:36]
  wire  _GEN_5260 = indexOnly ? _GEN_4228 : _GEN_4744; // @[dcache.scala 417:36]
  wire  _GEN_5261 = indexOnly ? _GEN_4229 : _GEN_4745; // @[dcache.scala 417:36]
  wire  _GEN_5262 = indexOnly ? _GEN_4230 : _GEN_4746; // @[dcache.scala 417:36]
  wire  _GEN_5263 = indexOnly ? _GEN_4231 : _GEN_4747; // @[dcache.scala 417:36]
  wire  _GEN_5264 = indexOnly ? _GEN_4232 : _GEN_4748; // @[dcache.scala 417:36]
  wire  _GEN_5265 = indexOnly ? _GEN_4233 : _GEN_4749; // @[dcache.scala 417:36]
  wire  _GEN_5266 = indexOnly ? _GEN_4234 : _GEN_4750; // @[dcache.scala 417:36]
  wire  _GEN_5267 = indexOnly ? _GEN_4235 : _GEN_4751; // @[dcache.scala 417:36]
  wire  _GEN_5268 = indexOnly ? _GEN_4236 : _GEN_4752; // @[dcache.scala 417:36]
  wire  _GEN_5269 = indexOnly ? _GEN_4237 : _GEN_4753; // @[dcache.scala 417:36]
  wire  _GEN_5270 = indexOnly ? _GEN_4238 : _GEN_4754; // @[dcache.scala 417:36]
  wire  _GEN_5271 = indexOnly ? _GEN_4239 : _GEN_4755; // @[dcache.scala 417:36]
  wire  _GEN_5272 = indexOnly ? _GEN_4240 : _GEN_4756; // @[dcache.scala 417:36]
  wire  _GEN_5273 = indexOnly ? _GEN_4241 : _GEN_4757; // @[dcache.scala 417:36]
  wire  _GEN_5274 = indexOnly ? _GEN_4242 : _GEN_4758; // @[dcache.scala 417:36]
  wire  _GEN_5275 = indexOnly ? _GEN_4243 : _GEN_4759; // @[dcache.scala 417:36]
  wire  _GEN_5276 = indexOnly ? _GEN_4244 : _GEN_4760; // @[dcache.scala 417:36]
  wire  _GEN_5277 = indexOnly ? _GEN_4245 : _GEN_4761; // @[dcache.scala 417:36]
  wire  _GEN_5278 = indexOnly ? _GEN_4246 : _GEN_4762; // @[dcache.scala 417:36]
  wire  _GEN_5279 = indexOnly ? _GEN_4247 : _GEN_4763; // @[dcache.scala 417:36]
  wire  _GEN_5280 = indexOnly ? _GEN_4248 : _GEN_4764; // @[dcache.scala 417:36]
  wire  _GEN_5281 = indexOnly ? _GEN_4249 : _GEN_4765; // @[dcache.scala 417:36]
  wire  _GEN_5282 = indexOnly ? _GEN_4250 : _GEN_4766; // @[dcache.scala 417:36]
  wire  _GEN_5283 = indexOnly ? _GEN_4251 : _GEN_4767; // @[dcache.scala 417:36]
  wire  _GEN_5284 = indexOnly ? _GEN_4252 : _GEN_4768; // @[dcache.scala 417:36]
  wire  _GEN_5285 = indexOnly ? _GEN_4253 : _GEN_4769; // @[dcache.scala 417:36]
  wire  _GEN_5286 = indexOnly ? _GEN_4254 : _GEN_4770; // @[dcache.scala 417:36]
  wire  _GEN_5287 = indexOnly ? _GEN_4255 : _GEN_4771; // @[dcache.scala 417:36]
  wire  _GEN_5288 = indexOnly ? _GEN_4256 : _GEN_4772; // @[dcache.scala 417:36]
  wire  _GEN_5289 = indexOnly ? _GEN_4257 : _GEN_4773; // @[dcache.scala 417:36]
  wire  _GEN_5290 = indexOnly ? _GEN_4258 : _GEN_4774; // @[dcache.scala 417:36]
  wire  _GEN_5291 = indexOnly ? _GEN_4259 : _GEN_4775; // @[dcache.scala 417:36]
  wire  _GEN_5292 = indexOnly ? _GEN_4260 : _GEN_4776; // @[dcache.scala 417:36]
  wire  _GEN_5293 = indexOnly ? _GEN_4261 : _GEN_4777; // @[dcache.scala 417:36]
  wire  _GEN_5294 = indexOnly ? _GEN_4262 : _GEN_4778; // @[dcache.scala 417:36]
  wire  _GEN_5295 = indexOnly ? _GEN_4263 : _GEN_4779; // @[dcache.scala 417:36]
  wire  _GEN_5296 = indexOnly ? _GEN_4264 : _GEN_4780; // @[dcache.scala 417:36]
  wire  _GEN_5297 = indexOnly ? _GEN_4265 : _GEN_4781; // @[dcache.scala 417:36]
  wire  _GEN_5298 = indexOnly ? _GEN_4266 : _GEN_4782; // @[dcache.scala 417:36]
  wire  _GEN_5299 = indexOnly ? _GEN_4267 : _GEN_4783; // @[dcache.scala 417:36]
  wire  _GEN_5300 = indexOnly ? _GEN_4268 : _GEN_4784; // @[dcache.scala 417:36]
  wire  _GEN_5301 = indexOnly ? _GEN_4269 : _GEN_4785; // @[dcache.scala 417:36]
  wire  _GEN_5302 = indexOnly ? _GEN_4270 : _GEN_4786; // @[dcache.scala 417:36]
  wire  _GEN_5303 = indexOnly ? _GEN_4271 : _GEN_4787; // @[dcache.scala 417:36]
  wire  _GEN_5304 = indexOnly ? _GEN_4272 : _GEN_4788; // @[dcache.scala 417:36]
  wire  _GEN_5305 = indexOnly ? _GEN_4273 : _GEN_4789; // @[dcache.scala 417:36]
  wire  _GEN_5306 = indexOnly ? _GEN_4274 : _GEN_4790; // @[dcache.scala 417:36]
  wire  _GEN_5307 = indexOnly ? _GEN_4275 : _GEN_4791; // @[dcache.scala 417:36]
  wire  _GEN_5308 = indexOnly ? _GEN_4276 : _GEN_4792; // @[dcache.scala 417:36]
  wire  _GEN_5309 = indexOnly ? _GEN_4277 : _GEN_4793; // @[dcache.scala 417:36]
  wire  _GEN_5310 = indexOnly ? _GEN_4278 : _GEN_4794; // @[dcache.scala 417:36]
  wire  _GEN_5311 = indexOnly ? _GEN_4279 : _GEN_4795; // @[dcache.scala 417:36]
  wire  _GEN_5312 = indexOnly ? _GEN_4280 : _GEN_4796; // @[dcache.scala 417:36]
  wire  _GEN_5313 = indexOnly ? _GEN_4281 : _GEN_4797; // @[dcache.scala 417:36]
  wire  _GEN_5314 = indexOnly ? _GEN_4282 : _GEN_4798; // @[dcache.scala 417:36]
  wire  _GEN_5315 = indexOnly ? _GEN_4283 : _GEN_4799; // @[dcache.scala 417:36]
  wire  _GEN_5316 = indexOnly ? _GEN_4284 : _GEN_4800; // @[dcache.scala 417:36]
  wire  _GEN_5317 = indexOnly ? _GEN_4285 : _GEN_4801; // @[dcache.scala 417:36]
  wire  _GEN_5318 = indexOnly ? _GEN_4286 : _GEN_4802; // @[dcache.scala 417:36]
  wire  _GEN_5319 = indexOnly ? _GEN_4287 : _GEN_4803; // @[dcache.scala 417:36]
  wire  _GEN_5320 = indexOnly ? _GEN_4288 : _GEN_4804; // @[dcache.scala 417:36]
  wire  _GEN_5321 = indexOnly ? _GEN_4289 : _GEN_4805; // @[dcache.scala 417:36]
  wire  _GEN_5322 = indexOnly ? _GEN_4290 : _GEN_4806; // @[dcache.scala 417:36]
  wire  _GEN_5323 = indexOnly ? _GEN_4291 : _GEN_4807; // @[dcache.scala 417:36]
  wire  _GEN_5324 = indexOnly ? _GEN_4292 : _GEN_4808; // @[dcache.scala 417:36]
  wire  _GEN_5325 = indexOnly ? _GEN_4293 : _GEN_4809; // @[dcache.scala 417:36]
  wire  _GEN_5326 = indexOnly ? _GEN_4294 : _GEN_4810; // @[dcache.scala 417:36]
  wire  _GEN_5327 = indexOnly ? _GEN_4295 : _GEN_4811; // @[dcache.scala 417:36]
  wire  _GEN_5328 = indexOnly ? _GEN_4296 : _GEN_4812; // @[dcache.scala 417:36]
  wire  _GEN_5329 = indexOnly ? _GEN_4297 : _GEN_4813; // @[dcache.scala 417:36]
  wire  _GEN_5330 = indexOnly ? _GEN_4298 : _GEN_4814; // @[dcache.scala 417:36]
  wire  _GEN_5331 = indexOnly ? _GEN_4299 : _GEN_4815; // @[dcache.scala 417:36]
  wire  _GEN_5332 = indexOnly ? _GEN_4300 : _GEN_4816; // @[dcache.scala 417:36]
  wire  _GEN_5333 = indexOnly ? _GEN_4301 : _GEN_4817; // @[dcache.scala 417:36]
  wire  _GEN_5334 = indexOnly ? _GEN_4302 : _GEN_4818; // @[dcache.scala 417:36]
  wire  _GEN_5335 = indexOnly ? _GEN_4303 : _GEN_4819; // @[dcache.scala 417:36]
  wire  _GEN_5336 = indexOnly ? _GEN_4304 : _GEN_4820; // @[dcache.scala 417:36]
  wire  _GEN_5337 = indexOnly ? _GEN_4305 : _GEN_4821; // @[dcache.scala 417:36]
  wire  _GEN_5338 = indexOnly ? _GEN_4306 : _GEN_4822; // @[dcache.scala 417:36]
  wire  _GEN_5339 = indexOnly ? _GEN_4307 : _GEN_4823; // @[dcache.scala 417:36]
  wire  _GEN_5340 = indexOnly ? _GEN_4308 : _GEN_4824; // @[dcache.scala 417:36]
  wire  _GEN_5341 = indexOnly ? _GEN_4309 : _GEN_4825; // @[dcache.scala 417:36]
  wire  _GEN_5342 = indexOnly ? _GEN_4310 : _GEN_4826; // @[dcache.scala 417:36]
  wire  _GEN_5343 = indexOnly ? _GEN_4311 : _GEN_4827; // @[dcache.scala 417:36]
  wire  _GEN_5344 = indexOnly ? _GEN_4312 : _GEN_4828; // @[dcache.scala 417:36]
  wire  _GEN_5345 = indexOnly ? _GEN_4313 : _GEN_4829; // @[dcache.scala 417:36]
  wire  _GEN_5346 = indexOnly ? _GEN_4314 : _GEN_4830; // @[dcache.scala 417:36]
  wire  _GEN_5347 = indexOnly ? _GEN_4315 : _GEN_4831; // @[dcache.scala 417:36]
  wire  _GEN_5348 = indexOnly ? _GEN_4316 : _GEN_4832; // @[dcache.scala 417:36]
  wire  _GEN_5349 = indexOnly ? _GEN_4317 : _GEN_4833; // @[dcache.scala 417:36]
  wire  _GEN_5350 = indexOnly ? _GEN_4318 : _GEN_4834; // @[dcache.scala 417:36]
  wire  _GEN_5351 = indexOnly ? _GEN_4319 : _GEN_4835; // @[dcache.scala 417:36]
  wire  _GEN_5352 = indexOnly ? _GEN_4320 : _GEN_4836; // @[dcache.scala 417:36]
  wire  _GEN_5353 = indexOnly ? _GEN_4321 : _GEN_4837; // @[dcache.scala 417:36]
  wire  _GEN_5354 = indexOnly ? _GEN_4322 : _GEN_4838; // @[dcache.scala 417:36]
  wire  _GEN_5355 = indexOnly ? _GEN_4323 : _GEN_4839; // @[dcache.scala 417:36]
  wire  _GEN_5356 = indexOnly ? _GEN_4324 : _GEN_4840; // @[dcache.scala 417:36]
  wire  _GEN_5357 = indexOnly ? _GEN_4325 : _GEN_4841; // @[dcache.scala 417:36]
  wire  _GEN_5358 = indexOnly ? _GEN_4326 : _GEN_4842; // @[dcache.scala 417:36]
  wire  _GEN_5359 = indexOnly ? _GEN_4327 : _GEN_4843; // @[dcache.scala 417:36]
  wire  _GEN_5360 = indexOnly ? _GEN_4328 : _GEN_4844; // @[dcache.scala 417:36]
  wire  _GEN_5361 = indexOnly ? _GEN_4329 : _GEN_4845; // @[dcache.scala 417:36]
  wire  _GEN_5362 = indexOnly ? _GEN_4330 : _GEN_4846; // @[dcache.scala 417:36]
  wire  _GEN_5363 = indexOnly ? _GEN_4331 : _GEN_4847; // @[dcache.scala 417:36]
  wire  _GEN_5364 = indexOnly ? _GEN_4332 : _GEN_4848; // @[dcache.scala 417:36]
  wire  _GEN_5365 = indexOnly ? _GEN_4333 : _GEN_4849; // @[dcache.scala 417:36]
  wire  _GEN_5366 = indexOnly ? _GEN_4334 : _GEN_4850; // @[dcache.scala 417:36]
  wire  _GEN_5367 = indexOnly ? _GEN_4335 : _GEN_4851; // @[dcache.scala 417:36]
  wire  _GEN_5368 = indexOnly ? _GEN_4336 : _GEN_4852; // @[dcache.scala 417:36]
  wire  _GEN_5369 = indexOnly ? _GEN_4337 : _GEN_4853; // @[dcache.scala 417:36]
  wire  _GEN_5370 = indexOnly ? _GEN_4338 : _GEN_4854; // @[dcache.scala 417:36]
  wire  _GEN_5371 = indexOnly ? _GEN_4339 : _GEN_4855; // @[dcache.scala 417:36]
  wire  _GEN_5372 = indexOnly ? _GEN_4340 : _GEN_4856; // @[dcache.scala 417:36]
  wire  _GEN_5373 = indexOnly ? _GEN_4341 : _GEN_4857; // @[dcache.scala 417:36]
  wire  _GEN_5374 = indexOnly ? _GEN_4342 : _GEN_4858; // @[dcache.scala 417:36]
  wire  _GEN_5375 = indexOnly ? _GEN_4343 : _GEN_4859; // @[dcache.scala 417:36]
  wire  _GEN_5376 = indexOnly ? _GEN_4344 : _GEN_4860; // @[dcache.scala 417:36]
  wire  _GEN_5377 = indexOnly ? _GEN_4345 : _GEN_4861; // @[dcache.scala 417:36]
  wire  _GEN_5378 = indexOnly ? _GEN_4346 : _GEN_4862; // @[dcache.scala 417:36]
  wire  _GEN_5379 = indexOnly ? _GEN_4347 : _GEN_4863; // @[dcache.scala 417:36]
  wire  _GEN_5380 = indexOnly ? _GEN_4348 : _GEN_4864; // @[dcache.scala 417:36]
  wire  _GEN_5381 = indexOnly ? _GEN_4349 : _GEN_4865; // @[dcache.scala 417:36]
  wire  _GEN_5382 = indexOnly ? _GEN_4350 : _GEN_4866; // @[dcache.scala 417:36]
  wire  _GEN_5383 = indexOnly ? _GEN_4351 : _GEN_4867; // @[dcache.scala 417:36]
  wire  _GEN_5384 = indexOnly ? _GEN_4352 : _GEN_4868; // @[dcache.scala 417:36]
  wire  _GEN_5385 = indexOnly ? _GEN_4353 : _GEN_4869; // @[dcache.scala 417:36]
  wire  _GEN_5386 = indexOnly ? _GEN_4354 : _GEN_4870; // @[dcache.scala 417:36]
  wire  _GEN_5387 = indexOnly ? _GEN_4355 : _GEN_4871; // @[dcache.scala 417:36]
  wire  _GEN_5388 = indexOnly ? _GEN_4356 : _GEN_4872; // @[dcache.scala 417:36]
  wire  _GEN_5389 = indexOnly ? _GEN_4357 : _GEN_4873; // @[dcache.scala 417:36]
  wire  _GEN_5390 = indexOnly ? _GEN_4358 : _GEN_4874; // @[dcache.scala 417:36]
  wire  _GEN_5391 = indexOnly ? _GEN_4359 : _GEN_4875; // @[dcache.scala 417:36]
  wire  _GEN_5392 = indexOnly ? _GEN_4360 : _GEN_4876; // @[dcache.scala 417:36]
  wire  _GEN_5393 = indexOnly ? _GEN_4361 : _GEN_4877; // @[dcache.scala 417:36]
  wire  _GEN_5394 = indexOnly ? _GEN_4362 : _GEN_4878; // @[dcache.scala 417:36]
  wire  _GEN_5395 = indexOnly ? _GEN_4363 : _GEN_4879; // @[dcache.scala 417:36]
  wire  _GEN_5396 = indexOnly ? _GEN_4364 : _GEN_4880; // @[dcache.scala 417:36]
  wire  _GEN_5397 = indexOnly ? _GEN_4365 : _GEN_4881; // @[dcache.scala 417:36]
  wire  _GEN_5398 = indexOnly ? _GEN_4366 : _GEN_4882; // @[dcache.scala 417:36]
  wire [20:0] _GEN_5399 = invalidate ? _GEN_4883 : _GEN_3335; // @[dcache.scala 416:33]
  wire [20:0] _GEN_5400 = invalidate ? _GEN_4884 : _GEN_3336; // @[dcache.scala 416:33]
  wire  _GEN_5401 = invalidate ? _GEN_4885 : _GEN_3337; // @[dcache.scala 416:33]
  wire  _GEN_5402 = invalidate ? _GEN_4886 : _GEN_3338; // @[dcache.scala 416:33]
  wire  _GEN_5403 = invalidate ? _GEN_4887 : _GEN_3339; // @[dcache.scala 416:33]
  wire  _GEN_5404 = invalidate ? _GEN_4888 : _GEN_3340; // @[dcache.scala 416:33]
  wire  _GEN_5405 = invalidate ? _GEN_4889 : _GEN_3341; // @[dcache.scala 416:33]
  wire  _GEN_5406 = invalidate ? _GEN_4890 : _GEN_3342; // @[dcache.scala 416:33]
  wire  _GEN_5407 = invalidate ? _GEN_4891 : _GEN_3343; // @[dcache.scala 416:33]
  wire  _GEN_5408 = invalidate ? _GEN_4892 : _GEN_3344; // @[dcache.scala 416:33]
  wire  _GEN_5409 = invalidate ? _GEN_4893 : _GEN_3345; // @[dcache.scala 416:33]
  wire  _GEN_5410 = invalidate ? _GEN_4894 : _GEN_3346; // @[dcache.scala 416:33]
  wire  _GEN_5411 = invalidate ? _GEN_4895 : _GEN_3347; // @[dcache.scala 416:33]
  wire  _GEN_5412 = invalidate ? _GEN_4896 : _GEN_3348; // @[dcache.scala 416:33]
  wire  _GEN_5413 = invalidate ? _GEN_4897 : _GEN_3349; // @[dcache.scala 416:33]
  wire  _GEN_5414 = invalidate ? _GEN_4898 : _GEN_3350; // @[dcache.scala 416:33]
  wire  _GEN_5415 = invalidate ? _GEN_4899 : _GEN_3351; // @[dcache.scala 416:33]
  wire  _GEN_5416 = invalidate ? _GEN_4900 : _GEN_3352; // @[dcache.scala 416:33]
  wire  _GEN_5417 = invalidate ? _GEN_4901 : _GEN_3353; // @[dcache.scala 416:33]
  wire  _GEN_5418 = invalidate ? _GEN_4902 : _GEN_3354; // @[dcache.scala 416:33]
  wire  _GEN_5419 = invalidate ? _GEN_4903 : _GEN_3355; // @[dcache.scala 416:33]
  wire  _GEN_5420 = invalidate ? _GEN_4904 : _GEN_3356; // @[dcache.scala 416:33]
  wire  _GEN_5421 = invalidate ? _GEN_4905 : _GEN_3357; // @[dcache.scala 416:33]
  wire  _GEN_5422 = invalidate ? _GEN_4906 : _GEN_3358; // @[dcache.scala 416:33]
  wire  _GEN_5423 = invalidate ? _GEN_4907 : _GEN_3359; // @[dcache.scala 416:33]
  wire  _GEN_5424 = invalidate ? _GEN_4908 : _GEN_3360; // @[dcache.scala 416:33]
  wire  _GEN_5425 = invalidate ? _GEN_4909 : _GEN_3361; // @[dcache.scala 416:33]
  wire  _GEN_5426 = invalidate ? _GEN_4910 : _GEN_3362; // @[dcache.scala 416:33]
  wire  _GEN_5427 = invalidate ? _GEN_4911 : _GEN_3363; // @[dcache.scala 416:33]
  wire  _GEN_5428 = invalidate ? _GEN_4912 : _GEN_3364; // @[dcache.scala 416:33]
  wire  _GEN_5429 = invalidate ? _GEN_4913 : _GEN_3365; // @[dcache.scala 416:33]
  wire  _GEN_5430 = invalidate ? _GEN_4914 : _GEN_3366; // @[dcache.scala 416:33]
  wire  _GEN_5431 = invalidate ? _GEN_4915 : _GEN_3367; // @[dcache.scala 416:33]
  wire  _GEN_5432 = invalidate ? _GEN_4916 : _GEN_3368; // @[dcache.scala 416:33]
  wire  _GEN_5433 = invalidate ? _GEN_4917 : _GEN_3369; // @[dcache.scala 416:33]
  wire  _GEN_5434 = invalidate ? _GEN_4918 : _GEN_3370; // @[dcache.scala 416:33]
  wire  _GEN_5435 = invalidate ? _GEN_4919 : _GEN_3371; // @[dcache.scala 416:33]
  wire  _GEN_5436 = invalidate ? _GEN_4920 : _GEN_3372; // @[dcache.scala 416:33]
  wire  _GEN_5437 = invalidate ? _GEN_4921 : _GEN_3373; // @[dcache.scala 416:33]
  wire  _GEN_5438 = invalidate ? _GEN_4922 : _GEN_3374; // @[dcache.scala 416:33]
  wire  _GEN_5439 = invalidate ? _GEN_4923 : _GEN_3375; // @[dcache.scala 416:33]
  wire  _GEN_5440 = invalidate ? _GEN_4924 : _GEN_3376; // @[dcache.scala 416:33]
  wire  _GEN_5441 = invalidate ? _GEN_4925 : _GEN_3377; // @[dcache.scala 416:33]
  wire  _GEN_5442 = invalidate ? _GEN_4926 : _GEN_3378; // @[dcache.scala 416:33]
  wire  _GEN_5443 = invalidate ? _GEN_4927 : _GEN_3379; // @[dcache.scala 416:33]
  wire  _GEN_5444 = invalidate ? _GEN_4928 : _GEN_3380; // @[dcache.scala 416:33]
  wire  _GEN_5445 = invalidate ? _GEN_4929 : _GEN_3381; // @[dcache.scala 416:33]
  wire  _GEN_5446 = invalidate ? _GEN_4930 : _GEN_3382; // @[dcache.scala 416:33]
  wire  _GEN_5447 = invalidate ? _GEN_4931 : _GEN_3383; // @[dcache.scala 416:33]
  wire  _GEN_5448 = invalidate ? _GEN_4932 : _GEN_3384; // @[dcache.scala 416:33]
  wire  _GEN_5449 = invalidate ? _GEN_4933 : _GEN_3385; // @[dcache.scala 416:33]
  wire  _GEN_5450 = invalidate ? _GEN_4934 : _GEN_3386; // @[dcache.scala 416:33]
  wire  _GEN_5451 = invalidate ? _GEN_4935 : _GEN_3387; // @[dcache.scala 416:33]
  wire  _GEN_5452 = invalidate ? _GEN_4936 : _GEN_3388; // @[dcache.scala 416:33]
  wire  _GEN_5453 = invalidate ? _GEN_4937 : _GEN_3389; // @[dcache.scala 416:33]
  wire  _GEN_5454 = invalidate ? _GEN_4938 : _GEN_3390; // @[dcache.scala 416:33]
  wire  _GEN_5455 = invalidate ? _GEN_4939 : _GEN_3391; // @[dcache.scala 416:33]
  wire  _GEN_5456 = invalidate ? _GEN_4940 : _GEN_3392; // @[dcache.scala 416:33]
  wire  _GEN_5457 = invalidate ? _GEN_4941 : _GEN_3393; // @[dcache.scala 416:33]
  wire  _GEN_5458 = invalidate ? _GEN_4942 : _GEN_3394; // @[dcache.scala 416:33]
  wire  _GEN_5459 = invalidate ? _GEN_4943 : _GEN_3395; // @[dcache.scala 416:33]
  wire  _GEN_5460 = invalidate ? _GEN_4944 : _GEN_3396; // @[dcache.scala 416:33]
  wire  _GEN_5461 = invalidate ? _GEN_4945 : _GEN_3397; // @[dcache.scala 416:33]
  wire  _GEN_5462 = invalidate ? _GEN_4946 : _GEN_3398; // @[dcache.scala 416:33]
  wire  _GEN_5463 = invalidate ? _GEN_4947 : _GEN_3399; // @[dcache.scala 416:33]
  wire  _GEN_5464 = invalidate ? _GEN_4948 : _GEN_3400; // @[dcache.scala 416:33]
  wire  _GEN_5465 = invalidate ? _GEN_4949 : _GEN_3401; // @[dcache.scala 416:33]
  wire  _GEN_5466 = invalidate ? _GEN_4950 : _GEN_3402; // @[dcache.scala 416:33]
  wire  _GEN_5467 = invalidate ? _GEN_4951 : _GEN_3403; // @[dcache.scala 416:33]
  wire  _GEN_5468 = invalidate ? _GEN_4952 : _GEN_3404; // @[dcache.scala 416:33]
  wire  _GEN_5469 = invalidate ? _GEN_4953 : _GEN_3405; // @[dcache.scala 416:33]
  wire  _GEN_5470 = invalidate ? _GEN_4954 : _GEN_3406; // @[dcache.scala 416:33]
  wire  _GEN_5471 = invalidate ? _GEN_4955 : _GEN_3407; // @[dcache.scala 416:33]
  wire  _GEN_5472 = invalidate ? _GEN_4956 : _GEN_3408; // @[dcache.scala 416:33]
  wire  _GEN_5473 = invalidate ? _GEN_4957 : _GEN_3409; // @[dcache.scala 416:33]
  wire  _GEN_5474 = invalidate ? _GEN_4958 : _GEN_3410; // @[dcache.scala 416:33]
  wire  _GEN_5475 = invalidate ? _GEN_4959 : _GEN_3411; // @[dcache.scala 416:33]
  wire  _GEN_5476 = invalidate ? _GEN_4960 : _GEN_3412; // @[dcache.scala 416:33]
  wire  _GEN_5477 = invalidate ? _GEN_4961 : _GEN_3413; // @[dcache.scala 416:33]
  wire  _GEN_5478 = invalidate ? _GEN_4962 : _GEN_3414; // @[dcache.scala 416:33]
  wire  _GEN_5479 = invalidate ? _GEN_4963 : _GEN_3415; // @[dcache.scala 416:33]
  wire  _GEN_5480 = invalidate ? _GEN_4964 : _GEN_3416; // @[dcache.scala 416:33]
  wire  _GEN_5481 = invalidate ? _GEN_4965 : _GEN_3417; // @[dcache.scala 416:33]
  wire  _GEN_5482 = invalidate ? _GEN_4966 : _GEN_3418; // @[dcache.scala 416:33]
  wire  _GEN_5483 = invalidate ? _GEN_4967 : _GEN_3419; // @[dcache.scala 416:33]
  wire  _GEN_5484 = invalidate ? _GEN_4968 : _GEN_3420; // @[dcache.scala 416:33]
  wire  _GEN_5485 = invalidate ? _GEN_4969 : _GEN_3421; // @[dcache.scala 416:33]
  wire  _GEN_5486 = invalidate ? _GEN_4970 : _GEN_3422; // @[dcache.scala 416:33]
  wire  _GEN_5487 = invalidate ? _GEN_4971 : _GEN_3423; // @[dcache.scala 416:33]
  wire  _GEN_5488 = invalidate ? _GEN_4972 : _GEN_3424; // @[dcache.scala 416:33]
  wire  _GEN_5489 = invalidate ? _GEN_4973 : _GEN_3425; // @[dcache.scala 416:33]
  wire  _GEN_5490 = invalidate ? _GEN_4974 : _GEN_3426; // @[dcache.scala 416:33]
  wire  _GEN_5491 = invalidate ? _GEN_4975 : _GEN_3427; // @[dcache.scala 416:33]
  wire  _GEN_5492 = invalidate ? _GEN_4976 : _GEN_3428; // @[dcache.scala 416:33]
  wire  _GEN_5493 = invalidate ? _GEN_4977 : _GEN_3429; // @[dcache.scala 416:33]
  wire  _GEN_5494 = invalidate ? _GEN_4978 : _GEN_3430; // @[dcache.scala 416:33]
  wire  _GEN_5495 = invalidate ? _GEN_4979 : _GEN_3431; // @[dcache.scala 416:33]
  wire  _GEN_5496 = invalidate ? _GEN_4980 : _GEN_3432; // @[dcache.scala 416:33]
  wire  _GEN_5497 = invalidate ? _GEN_4981 : _GEN_3433; // @[dcache.scala 416:33]
  wire  _GEN_5498 = invalidate ? _GEN_4982 : _GEN_3434; // @[dcache.scala 416:33]
  wire  _GEN_5499 = invalidate ? _GEN_4983 : _GEN_3435; // @[dcache.scala 416:33]
  wire  _GEN_5500 = invalidate ? _GEN_4984 : _GEN_3436; // @[dcache.scala 416:33]
  wire  _GEN_5501 = invalidate ? _GEN_4985 : _GEN_3437; // @[dcache.scala 416:33]
  wire  _GEN_5502 = invalidate ? _GEN_4986 : _GEN_3438; // @[dcache.scala 416:33]
  wire  _GEN_5503 = invalidate ? _GEN_4987 : _GEN_3439; // @[dcache.scala 416:33]
  wire  _GEN_5504 = invalidate ? _GEN_4988 : _GEN_3440; // @[dcache.scala 416:33]
  wire  _GEN_5505 = invalidate ? _GEN_4989 : _GEN_3441; // @[dcache.scala 416:33]
  wire  _GEN_5506 = invalidate ? _GEN_4990 : _GEN_3442; // @[dcache.scala 416:33]
  wire  _GEN_5507 = invalidate ? _GEN_4991 : _GEN_3443; // @[dcache.scala 416:33]
  wire  _GEN_5508 = invalidate ? _GEN_4992 : _GEN_3444; // @[dcache.scala 416:33]
  wire  _GEN_5509 = invalidate ? _GEN_4993 : _GEN_3445; // @[dcache.scala 416:33]
  wire  _GEN_5510 = invalidate ? _GEN_4994 : _GEN_3446; // @[dcache.scala 416:33]
  wire  _GEN_5511 = invalidate ? _GEN_4995 : _GEN_3447; // @[dcache.scala 416:33]
  wire  _GEN_5512 = invalidate ? _GEN_4996 : _GEN_3448; // @[dcache.scala 416:33]
  wire  _GEN_5513 = invalidate ? _GEN_4997 : _GEN_3449; // @[dcache.scala 416:33]
  wire  _GEN_5514 = invalidate ? _GEN_4998 : _GEN_3450; // @[dcache.scala 416:33]
  wire  _GEN_5515 = invalidate ? _GEN_4999 : _GEN_3451; // @[dcache.scala 416:33]
  wire  _GEN_5516 = invalidate ? _GEN_5000 : _GEN_3452; // @[dcache.scala 416:33]
  wire  _GEN_5517 = invalidate ? _GEN_5001 : _GEN_3453; // @[dcache.scala 416:33]
  wire  _GEN_5518 = invalidate ? _GEN_5002 : _GEN_3454; // @[dcache.scala 416:33]
  wire  _GEN_5519 = invalidate ? _GEN_5003 : _GEN_3455; // @[dcache.scala 416:33]
  wire  _GEN_5520 = invalidate ? _GEN_5004 : _GEN_3456; // @[dcache.scala 416:33]
  wire  _GEN_5521 = invalidate ? _GEN_5005 : _GEN_3457; // @[dcache.scala 416:33]
  wire  _GEN_5522 = invalidate ? _GEN_5006 : _GEN_3458; // @[dcache.scala 416:33]
  wire  _GEN_5523 = invalidate ? _GEN_5007 : _GEN_3459; // @[dcache.scala 416:33]
  wire  _GEN_5524 = invalidate ? _GEN_5008 : _GEN_3460; // @[dcache.scala 416:33]
  wire  _GEN_5525 = invalidate ? _GEN_5009 : _GEN_3461; // @[dcache.scala 416:33]
  wire  _GEN_5526 = invalidate ? _GEN_5010 : _GEN_3462; // @[dcache.scala 416:33]
  wire  _GEN_5527 = invalidate ? _GEN_5011 : _GEN_3463; // @[dcache.scala 416:33]
  wire  _GEN_5528 = invalidate ? _GEN_5012 : _GEN_3464; // @[dcache.scala 416:33]
  wire  _GEN_5529 = invalidate ? _GEN_5013 : _GEN_3465; // @[dcache.scala 416:33]
  wire  _GEN_5530 = invalidate ? _GEN_5014 : _GEN_3466; // @[dcache.scala 416:33]
  wire  _GEN_5531 = invalidate ? _GEN_5015 : _GEN_3467; // @[dcache.scala 416:33]
  wire  _GEN_5532 = invalidate ? _GEN_5016 : _GEN_3468; // @[dcache.scala 416:33]
  wire  _GEN_5533 = invalidate ? _GEN_5017 : _GEN_3469; // @[dcache.scala 416:33]
  wire  _GEN_5534 = invalidate ? _GEN_5018 : _GEN_3470; // @[dcache.scala 416:33]
  wire  _GEN_5535 = invalidate ? _GEN_5019 : _GEN_3471; // @[dcache.scala 416:33]
  wire  _GEN_5536 = invalidate ? _GEN_5020 : _GEN_3472; // @[dcache.scala 416:33]
  wire  _GEN_5537 = invalidate ? _GEN_5021 : _GEN_3473; // @[dcache.scala 416:33]
  wire  _GEN_5538 = invalidate ? _GEN_5022 : _GEN_3474; // @[dcache.scala 416:33]
  wire  _GEN_5539 = invalidate ? _GEN_5023 : _GEN_3475; // @[dcache.scala 416:33]
  wire  _GEN_5540 = invalidate ? _GEN_5024 : _GEN_3476; // @[dcache.scala 416:33]
  wire  _GEN_5541 = invalidate ? _GEN_5025 : _GEN_3477; // @[dcache.scala 416:33]
  wire  _GEN_5542 = invalidate ? _GEN_5026 : _GEN_3478; // @[dcache.scala 416:33]
  wire  _GEN_5543 = invalidate ? _GEN_5027 : _GEN_3479; // @[dcache.scala 416:33]
  wire  _GEN_5544 = invalidate ? _GEN_5028 : _GEN_3480; // @[dcache.scala 416:33]
  wire  _GEN_5545 = invalidate ? _GEN_5029 : _GEN_3481; // @[dcache.scala 416:33]
  wire  _GEN_5546 = invalidate ? _GEN_5030 : _GEN_3482; // @[dcache.scala 416:33]
  wire  _GEN_5547 = invalidate ? _GEN_5031 : _GEN_3483; // @[dcache.scala 416:33]
  wire  _GEN_5548 = invalidate ? _GEN_5032 : _GEN_3484; // @[dcache.scala 416:33]
  wire  _GEN_5549 = invalidate ? _GEN_5033 : _GEN_3485; // @[dcache.scala 416:33]
  wire  _GEN_5550 = invalidate ? _GEN_5034 : _GEN_3486; // @[dcache.scala 416:33]
  wire  _GEN_5551 = invalidate ? _GEN_5035 : _GEN_3487; // @[dcache.scala 416:33]
  wire  _GEN_5552 = invalidate ? _GEN_5036 : _GEN_3488; // @[dcache.scala 416:33]
  wire  _GEN_5553 = invalidate ? _GEN_5037 : _GEN_3489; // @[dcache.scala 416:33]
  wire  _GEN_5554 = invalidate ? _GEN_5038 : _GEN_3490; // @[dcache.scala 416:33]
  wire  _GEN_5555 = invalidate ? _GEN_5039 : _GEN_3491; // @[dcache.scala 416:33]
  wire  _GEN_5556 = invalidate ? _GEN_5040 : _GEN_3492; // @[dcache.scala 416:33]
  wire  _GEN_5557 = invalidate ? _GEN_5041 : _GEN_3493; // @[dcache.scala 416:33]
  wire  _GEN_5558 = invalidate ? _GEN_5042 : _GEN_3494; // @[dcache.scala 416:33]
  wire  _GEN_5559 = invalidate ? _GEN_5043 : _GEN_3495; // @[dcache.scala 416:33]
  wire  _GEN_5560 = invalidate ? _GEN_5044 : _GEN_3496; // @[dcache.scala 416:33]
  wire  _GEN_5561 = invalidate ? _GEN_5045 : _GEN_3497; // @[dcache.scala 416:33]
  wire  _GEN_5562 = invalidate ? _GEN_5046 : _GEN_3498; // @[dcache.scala 416:33]
  wire  _GEN_5563 = invalidate ? _GEN_5047 : _GEN_3499; // @[dcache.scala 416:33]
  wire  _GEN_5564 = invalidate ? _GEN_5048 : _GEN_3500; // @[dcache.scala 416:33]
  wire  _GEN_5565 = invalidate ? _GEN_5049 : _GEN_3501; // @[dcache.scala 416:33]
  wire  _GEN_5566 = invalidate ? _GEN_5050 : _GEN_3502; // @[dcache.scala 416:33]
  wire  _GEN_5567 = invalidate ? _GEN_5051 : _GEN_3503; // @[dcache.scala 416:33]
  wire  _GEN_5568 = invalidate ? _GEN_5052 : _GEN_3504; // @[dcache.scala 416:33]
  wire  _GEN_5569 = invalidate ? _GEN_5053 : _GEN_3505; // @[dcache.scala 416:33]
  wire  _GEN_5570 = invalidate ? _GEN_5054 : _GEN_3506; // @[dcache.scala 416:33]
  wire  _GEN_5571 = invalidate ? _GEN_5055 : _GEN_3507; // @[dcache.scala 416:33]
  wire  _GEN_5572 = invalidate ? _GEN_5056 : _GEN_3508; // @[dcache.scala 416:33]
  wire  _GEN_5573 = invalidate ? _GEN_5057 : _GEN_3509; // @[dcache.scala 416:33]
  wire  _GEN_5574 = invalidate ? _GEN_5058 : _GEN_3510; // @[dcache.scala 416:33]
  wire  _GEN_5575 = invalidate ? _GEN_5059 : _GEN_3511; // @[dcache.scala 416:33]
  wire  _GEN_5576 = invalidate ? _GEN_5060 : _GEN_3512; // @[dcache.scala 416:33]
  wire  _GEN_5577 = invalidate ? _GEN_5061 : _GEN_3513; // @[dcache.scala 416:33]
  wire  _GEN_5578 = invalidate ? _GEN_5062 : _GEN_3514; // @[dcache.scala 416:33]
  wire  _GEN_5579 = invalidate ? _GEN_5063 : _GEN_3515; // @[dcache.scala 416:33]
  wire  _GEN_5580 = invalidate ? _GEN_5064 : _GEN_3516; // @[dcache.scala 416:33]
  wire  _GEN_5581 = invalidate ? _GEN_5065 : _GEN_3517; // @[dcache.scala 416:33]
  wire  _GEN_5582 = invalidate ? _GEN_5066 : _GEN_3518; // @[dcache.scala 416:33]
  wire  _GEN_5583 = invalidate ? _GEN_5067 : _GEN_3519; // @[dcache.scala 416:33]
  wire  _GEN_5584 = invalidate ? _GEN_5068 : _GEN_3520; // @[dcache.scala 416:33]
  wire  _GEN_5585 = invalidate ? _GEN_5069 : _GEN_3521; // @[dcache.scala 416:33]
  wire  _GEN_5586 = invalidate ? _GEN_5070 : _GEN_3522; // @[dcache.scala 416:33]
  wire  _GEN_5587 = invalidate ? _GEN_5071 : _GEN_3523; // @[dcache.scala 416:33]
  wire  _GEN_5588 = invalidate ? _GEN_5072 : _GEN_3524; // @[dcache.scala 416:33]
  wire  _GEN_5589 = invalidate ? _GEN_5073 : _GEN_3525; // @[dcache.scala 416:33]
  wire  _GEN_5590 = invalidate ? _GEN_5074 : _GEN_3526; // @[dcache.scala 416:33]
  wire  _GEN_5591 = invalidate ? _GEN_5075 : _GEN_3527; // @[dcache.scala 416:33]
  wire  _GEN_5592 = invalidate ? _GEN_5076 : _GEN_3528; // @[dcache.scala 416:33]
  wire  _GEN_5593 = invalidate ? _GEN_5077 : _GEN_3529; // @[dcache.scala 416:33]
  wire  _GEN_5594 = invalidate ? _GEN_5078 : _GEN_3530; // @[dcache.scala 416:33]
  wire  _GEN_5595 = invalidate ? _GEN_5079 : _GEN_3531; // @[dcache.scala 416:33]
  wire  _GEN_5596 = invalidate ? _GEN_5080 : _GEN_3532; // @[dcache.scala 416:33]
  wire  _GEN_5597 = invalidate ? _GEN_5081 : _GEN_3533; // @[dcache.scala 416:33]
  wire  _GEN_5598 = invalidate ? _GEN_5082 : _GEN_3534; // @[dcache.scala 416:33]
  wire  _GEN_5599 = invalidate ? _GEN_5083 : _GEN_3535; // @[dcache.scala 416:33]
  wire  _GEN_5600 = invalidate ? _GEN_5084 : _GEN_3536; // @[dcache.scala 416:33]
  wire  _GEN_5601 = invalidate ? _GEN_5085 : _GEN_3537; // @[dcache.scala 416:33]
  wire  _GEN_5602 = invalidate ? _GEN_5086 : _GEN_3538; // @[dcache.scala 416:33]
  wire  _GEN_5603 = invalidate ? _GEN_5087 : _GEN_3539; // @[dcache.scala 416:33]
  wire  _GEN_5604 = invalidate ? _GEN_5088 : _GEN_3540; // @[dcache.scala 416:33]
  wire  _GEN_5605 = invalidate ? _GEN_5089 : _GEN_3541; // @[dcache.scala 416:33]
  wire  _GEN_5606 = invalidate ? _GEN_5090 : _GEN_3542; // @[dcache.scala 416:33]
  wire  _GEN_5607 = invalidate ? _GEN_5091 : _GEN_3543; // @[dcache.scala 416:33]
  wire  _GEN_5608 = invalidate ? _GEN_5092 : _GEN_3544; // @[dcache.scala 416:33]
  wire  _GEN_5609 = invalidate ? _GEN_5093 : _GEN_3545; // @[dcache.scala 416:33]
  wire  _GEN_5610 = invalidate ? _GEN_5094 : _GEN_3546; // @[dcache.scala 416:33]
  wire  _GEN_5611 = invalidate ? _GEN_5095 : _GEN_3547; // @[dcache.scala 416:33]
  wire  _GEN_5612 = invalidate ? _GEN_5096 : _GEN_3548; // @[dcache.scala 416:33]
  wire  _GEN_5613 = invalidate ? _GEN_5097 : _GEN_3549; // @[dcache.scala 416:33]
  wire  _GEN_5614 = invalidate ? _GEN_5098 : _GEN_3550; // @[dcache.scala 416:33]
  wire  _GEN_5615 = invalidate ? _GEN_5099 : _GEN_3551; // @[dcache.scala 416:33]
  wire  _GEN_5616 = invalidate ? _GEN_5100 : _GEN_3552; // @[dcache.scala 416:33]
  wire  _GEN_5617 = invalidate ? _GEN_5101 : _GEN_3553; // @[dcache.scala 416:33]
  wire  _GEN_5618 = invalidate ? _GEN_5102 : _GEN_3554; // @[dcache.scala 416:33]
  wire  _GEN_5619 = invalidate ? _GEN_5103 : _GEN_3555; // @[dcache.scala 416:33]
  wire  _GEN_5620 = invalidate ? _GEN_5104 : _GEN_3556; // @[dcache.scala 416:33]
  wire  _GEN_5621 = invalidate ? _GEN_5105 : _GEN_3557; // @[dcache.scala 416:33]
  wire  _GEN_5622 = invalidate ? _GEN_5106 : _GEN_3558; // @[dcache.scala 416:33]
  wire  _GEN_5623 = invalidate ? _GEN_5107 : _GEN_3559; // @[dcache.scala 416:33]
  wire  _GEN_5624 = invalidate ? _GEN_5108 : _GEN_3560; // @[dcache.scala 416:33]
  wire  _GEN_5625 = invalidate ? _GEN_5109 : _GEN_3561; // @[dcache.scala 416:33]
  wire  _GEN_5626 = invalidate ? _GEN_5110 : _GEN_3562; // @[dcache.scala 416:33]
  wire  _GEN_5627 = invalidate ? _GEN_5111 : _GEN_3563; // @[dcache.scala 416:33]
  wire  _GEN_5628 = invalidate ? _GEN_5112 : _GEN_3564; // @[dcache.scala 416:33]
  wire  _GEN_5629 = invalidate ? _GEN_5113 : _GEN_3565; // @[dcache.scala 416:33]
  wire  _GEN_5630 = invalidate ? _GEN_5114 : _GEN_3566; // @[dcache.scala 416:33]
  wire  _GEN_5631 = invalidate ? _GEN_5115 : _GEN_3567; // @[dcache.scala 416:33]
  wire  _GEN_5632 = invalidate ? _GEN_5116 : _GEN_3568; // @[dcache.scala 416:33]
  wire  _GEN_5633 = invalidate ? _GEN_5117 : _GEN_3569; // @[dcache.scala 416:33]
  wire  _GEN_5634 = invalidate ? _GEN_5118 : _GEN_3570; // @[dcache.scala 416:33]
  wire  _GEN_5635 = invalidate ? _GEN_5119 : _GEN_3571; // @[dcache.scala 416:33]
  wire  _GEN_5636 = invalidate ? _GEN_5120 : _GEN_3572; // @[dcache.scala 416:33]
  wire  _GEN_5637 = invalidate ? _GEN_5121 : _GEN_3573; // @[dcache.scala 416:33]
  wire  _GEN_5638 = invalidate ? _GEN_5122 : _GEN_3574; // @[dcache.scala 416:33]
  wire  _GEN_5639 = invalidate ? _GEN_5123 : _GEN_3575; // @[dcache.scala 416:33]
  wire  _GEN_5640 = invalidate ? _GEN_5124 : _GEN_3576; // @[dcache.scala 416:33]
  wire  _GEN_5641 = invalidate ? _GEN_5125 : _GEN_3577; // @[dcache.scala 416:33]
  wire  _GEN_5642 = invalidate ? _GEN_5126 : _GEN_3578; // @[dcache.scala 416:33]
  wire  _GEN_5643 = invalidate ? _GEN_5127 : _GEN_3579; // @[dcache.scala 416:33]
  wire  _GEN_5644 = invalidate ? _GEN_5128 : _GEN_3580; // @[dcache.scala 416:33]
  wire  _GEN_5645 = invalidate ? _GEN_5129 : _GEN_3581; // @[dcache.scala 416:33]
  wire  _GEN_5646 = invalidate ? _GEN_5130 : _GEN_3582; // @[dcache.scala 416:33]
  wire  _GEN_5647 = invalidate ? _GEN_5131 : _GEN_3583; // @[dcache.scala 416:33]
  wire  _GEN_5648 = invalidate ? _GEN_5132 : _GEN_3584; // @[dcache.scala 416:33]
  wire  _GEN_5649 = invalidate ? _GEN_5133 : _GEN_3585; // @[dcache.scala 416:33]
  wire  _GEN_5650 = invalidate ? _GEN_5134 : _GEN_3586; // @[dcache.scala 416:33]
  wire  _GEN_5651 = invalidate ? _GEN_5135 : _GEN_3587; // @[dcache.scala 416:33]
  wire  _GEN_5652 = invalidate ? _GEN_5136 : _GEN_3588; // @[dcache.scala 416:33]
  wire  _GEN_5653 = invalidate ? _GEN_5137 : _GEN_3589; // @[dcache.scala 416:33]
  wire  _GEN_5654 = invalidate ? _GEN_5138 : _GEN_3590; // @[dcache.scala 416:33]
  wire  _GEN_5655 = invalidate ? _GEN_5139 : _GEN_3591; // @[dcache.scala 416:33]
  wire  _GEN_5656 = invalidate ? _GEN_5140 : _GEN_3592; // @[dcache.scala 416:33]
  wire  _GEN_5657 = invalidate ? _GEN_5141 : _GEN_3593; // @[dcache.scala 416:33]
  wire  _GEN_5658 = invalidate ? _GEN_5142 : _GEN_3594; // @[dcache.scala 416:33]
  wire  _GEN_5659 = invalidate ? _GEN_5143 : _GEN_3595; // @[dcache.scala 416:33]
  wire  _GEN_5660 = invalidate ? _GEN_5144 : _GEN_3596; // @[dcache.scala 416:33]
  wire  _GEN_5661 = invalidate ? _GEN_5145 : _GEN_3597; // @[dcache.scala 416:33]
  wire  _GEN_5662 = invalidate ? _GEN_5146 : _GEN_3598; // @[dcache.scala 416:33]
  wire  _GEN_5663 = invalidate ? _GEN_5147 : _GEN_3599; // @[dcache.scala 416:33]
  wire  _GEN_5664 = invalidate ? _GEN_5148 : _GEN_3600; // @[dcache.scala 416:33]
  wire  _GEN_5665 = invalidate ? _GEN_5149 : _GEN_3601; // @[dcache.scala 416:33]
  wire  _GEN_5666 = invalidate ? _GEN_5150 : _GEN_3602; // @[dcache.scala 416:33]
  wire  _GEN_5667 = invalidate ? _GEN_5151 : _GEN_3603; // @[dcache.scala 416:33]
  wire  _GEN_5668 = invalidate ? _GEN_5152 : _GEN_3604; // @[dcache.scala 416:33]
  wire  _GEN_5669 = invalidate ? _GEN_5153 : _GEN_3605; // @[dcache.scala 416:33]
  wire  _GEN_5670 = invalidate ? _GEN_5154 : _GEN_3606; // @[dcache.scala 416:33]
  wire  _GEN_5671 = invalidate ? _GEN_5155 : _GEN_3607; // @[dcache.scala 416:33]
  wire  _GEN_5672 = invalidate ? _GEN_5156 : _GEN_3608; // @[dcache.scala 416:33]
  wire  _GEN_5673 = invalidate ? _GEN_5157 : _GEN_3609; // @[dcache.scala 416:33]
  wire  _GEN_5674 = invalidate ? _GEN_5158 : _GEN_3610; // @[dcache.scala 416:33]
  wire  _GEN_5675 = invalidate ? _GEN_5159 : _GEN_3611; // @[dcache.scala 416:33]
  wire  _GEN_5676 = invalidate ? _GEN_5160 : _GEN_3612; // @[dcache.scala 416:33]
  wire  _GEN_5677 = invalidate ? _GEN_5161 : _GEN_3613; // @[dcache.scala 416:33]
  wire  _GEN_5678 = invalidate ? _GEN_5162 : _GEN_3614; // @[dcache.scala 416:33]
  wire  _GEN_5679 = invalidate ? _GEN_5163 : _GEN_3615; // @[dcache.scala 416:33]
  wire  _GEN_5680 = invalidate ? _GEN_5164 : _GEN_3616; // @[dcache.scala 416:33]
  wire  _GEN_5681 = invalidate ? _GEN_5165 : _GEN_3617; // @[dcache.scala 416:33]
  wire  _GEN_5682 = invalidate ? _GEN_5166 : _GEN_3618; // @[dcache.scala 416:33]
  wire  _GEN_5683 = invalidate ? _GEN_5167 : _GEN_3619; // @[dcache.scala 416:33]
  wire  _GEN_5684 = invalidate ? _GEN_5168 : _GEN_3620; // @[dcache.scala 416:33]
  wire  _GEN_5685 = invalidate ? _GEN_5169 : _GEN_3621; // @[dcache.scala 416:33]
  wire  _GEN_5686 = invalidate ? _GEN_5170 : _GEN_3622; // @[dcache.scala 416:33]
  wire  _GEN_5687 = invalidate ? _GEN_5171 : _GEN_3623; // @[dcache.scala 416:33]
  wire  _GEN_5688 = invalidate ? _GEN_5172 : _GEN_3624; // @[dcache.scala 416:33]
  wire  _GEN_5689 = invalidate ? _GEN_5173 : _GEN_3625; // @[dcache.scala 416:33]
  wire  _GEN_5690 = invalidate ? _GEN_5174 : _GEN_3626; // @[dcache.scala 416:33]
  wire  _GEN_5691 = invalidate ? _GEN_5175 : _GEN_3627; // @[dcache.scala 416:33]
  wire  _GEN_5692 = invalidate ? _GEN_5176 : _GEN_3628; // @[dcache.scala 416:33]
  wire  _GEN_5693 = invalidate ? _GEN_5177 : _GEN_3629; // @[dcache.scala 416:33]
  wire  _GEN_5694 = invalidate ? _GEN_5178 : _GEN_3630; // @[dcache.scala 416:33]
  wire  _GEN_5695 = invalidate ? _GEN_5179 : _GEN_3631; // @[dcache.scala 416:33]
  wire  _GEN_5696 = invalidate ? _GEN_5180 : _GEN_3632; // @[dcache.scala 416:33]
  wire  _GEN_5697 = invalidate ? _GEN_5181 : _GEN_3633; // @[dcache.scala 416:33]
  wire  _GEN_5698 = invalidate ? _GEN_5182 : _GEN_3634; // @[dcache.scala 416:33]
  wire  _GEN_5699 = invalidate ? _GEN_5183 : _GEN_3635; // @[dcache.scala 416:33]
  wire  _GEN_5700 = invalidate ? _GEN_5184 : _GEN_3636; // @[dcache.scala 416:33]
  wire  _GEN_5701 = invalidate ? _GEN_5185 : _GEN_3637; // @[dcache.scala 416:33]
  wire  _GEN_5702 = invalidate ? _GEN_5186 : _GEN_3638; // @[dcache.scala 416:33]
  wire  _GEN_5703 = invalidate ? _GEN_5187 : _GEN_3639; // @[dcache.scala 416:33]
  wire  _GEN_5704 = invalidate ? _GEN_5188 : _GEN_3640; // @[dcache.scala 416:33]
  wire  _GEN_5705 = invalidate ? _GEN_5189 : _GEN_3641; // @[dcache.scala 416:33]
  wire  _GEN_5706 = invalidate ? _GEN_5190 : _GEN_3642; // @[dcache.scala 416:33]
  wire  _GEN_5707 = invalidate ? _GEN_5191 : _GEN_3643; // @[dcache.scala 416:33]
  wire  _GEN_5708 = invalidate ? _GEN_5192 : _GEN_3644; // @[dcache.scala 416:33]
  wire  _GEN_5709 = invalidate ? _GEN_5193 : _GEN_3645; // @[dcache.scala 416:33]
  wire  _GEN_5710 = invalidate ? _GEN_5194 : _GEN_3646; // @[dcache.scala 416:33]
  wire  _GEN_5711 = invalidate ? _GEN_5195 : _GEN_3647; // @[dcache.scala 416:33]
  wire  _GEN_5712 = invalidate ? _GEN_5196 : _GEN_3648; // @[dcache.scala 416:33]
  wire  _GEN_5713 = invalidate ? _GEN_5197 : _GEN_3649; // @[dcache.scala 416:33]
  wire  _GEN_5714 = invalidate ? _GEN_5198 : _GEN_3650; // @[dcache.scala 416:33]
  wire  _GEN_5715 = invalidate ? _GEN_5199 : _GEN_3651; // @[dcache.scala 416:33]
  wire  _GEN_5716 = invalidate ? _GEN_5200 : _GEN_3652; // @[dcache.scala 416:33]
  wire  _GEN_5717 = invalidate ? _GEN_5201 : _GEN_3653; // @[dcache.scala 416:33]
  wire  _GEN_5718 = invalidate ? _GEN_5202 : _GEN_3654; // @[dcache.scala 416:33]
  wire  _GEN_5719 = invalidate ? _GEN_5203 : _GEN_3655; // @[dcache.scala 416:33]
  wire  _GEN_5720 = invalidate ? _GEN_5204 : _GEN_3656; // @[dcache.scala 416:33]
  wire  _GEN_5721 = invalidate ? _GEN_5205 : _GEN_3657; // @[dcache.scala 416:33]
  wire  _GEN_5722 = invalidate ? _GEN_5206 : _GEN_3658; // @[dcache.scala 416:33]
  wire  _GEN_5723 = invalidate ? _GEN_5207 : _GEN_3659; // @[dcache.scala 416:33]
  wire  _GEN_5724 = invalidate ? _GEN_5208 : _GEN_3660; // @[dcache.scala 416:33]
  wire  _GEN_5725 = invalidate ? _GEN_5209 : _GEN_3661; // @[dcache.scala 416:33]
  wire  _GEN_5726 = invalidate ? _GEN_5210 : _GEN_3662; // @[dcache.scala 416:33]
  wire  _GEN_5727 = invalidate ? _GEN_5211 : _GEN_3663; // @[dcache.scala 416:33]
  wire  _GEN_5728 = invalidate ? _GEN_5212 : _GEN_3664; // @[dcache.scala 416:33]
  wire  _GEN_5729 = invalidate ? _GEN_5213 : _GEN_3665; // @[dcache.scala 416:33]
  wire  _GEN_5730 = invalidate ? _GEN_5214 : _GEN_3666; // @[dcache.scala 416:33]
  wire  _GEN_5731 = invalidate ? _GEN_5215 : _GEN_3667; // @[dcache.scala 416:33]
  wire  _GEN_5732 = invalidate ? _GEN_5216 : _GEN_3668; // @[dcache.scala 416:33]
  wire  _GEN_5733 = invalidate ? _GEN_5217 : _GEN_3669; // @[dcache.scala 416:33]
  wire  _GEN_5734 = invalidate ? _GEN_5218 : _GEN_3670; // @[dcache.scala 416:33]
  wire  _GEN_5735 = invalidate ? _GEN_5219 : _GEN_3671; // @[dcache.scala 416:33]
  wire  _GEN_5736 = invalidate ? _GEN_5220 : _GEN_3672; // @[dcache.scala 416:33]
  wire  _GEN_5737 = invalidate ? _GEN_5221 : _GEN_3673; // @[dcache.scala 416:33]
  wire  _GEN_5738 = invalidate ? _GEN_5222 : _GEN_3674; // @[dcache.scala 416:33]
  wire  _GEN_5739 = invalidate ? _GEN_5223 : _GEN_3675; // @[dcache.scala 416:33]
  wire  _GEN_5740 = invalidate ? _GEN_5224 : _GEN_3676; // @[dcache.scala 416:33]
  wire  _GEN_5741 = invalidate ? _GEN_5225 : _GEN_3677; // @[dcache.scala 416:33]
  wire  _GEN_5742 = invalidate ? _GEN_5226 : _GEN_3678; // @[dcache.scala 416:33]
  wire  _GEN_5743 = invalidate ? _GEN_5227 : _GEN_3679; // @[dcache.scala 416:33]
  wire  _GEN_5744 = invalidate ? _GEN_5228 : _GEN_3680; // @[dcache.scala 416:33]
  wire  _GEN_5745 = invalidate ? _GEN_5229 : _GEN_3681; // @[dcache.scala 416:33]
  wire  _GEN_5746 = invalidate ? _GEN_5230 : _GEN_3682; // @[dcache.scala 416:33]
  wire  _GEN_5747 = invalidate ? _GEN_5231 : _GEN_3683; // @[dcache.scala 416:33]
  wire  _GEN_5748 = invalidate ? _GEN_5232 : _GEN_3684; // @[dcache.scala 416:33]
  wire  _GEN_5749 = invalidate ? _GEN_5233 : _GEN_3685; // @[dcache.scala 416:33]
  wire  _GEN_5750 = invalidate ? _GEN_5234 : _GEN_3686; // @[dcache.scala 416:33]
  wire  _GEN_5751 = invalidate ? _GEN_5235 : _GEN_3687; // @[dcache.scala 416:33]
  wire  _GEN_5752 = invalidate ? _GEN_5236 : _GEN_3688; // @[dcache.scala 416:33]
  wire  _GEN_5753 = invalidate ? _GEN_5237 : _GEN_3689; // @[dcache.scala 416:33]
  wire  _GEN_5754 = invalidate ? _GEN_5238 : _GEN_3690; // @[dcache.scala 416:33]
  wire  _GEN_5755 = invalidate ? _GEN_5239 : _GEN_3691; // @[dcache.scala 416:33]
  wire  _GEN_5756 = invalidate ? _GEN_5240 : _GEN_3692; // @[dcache.scala 416:33]
  wire  _GEN_5757 = invalidate ? _GEN_5241 : _GEN_3693; // @[dcache.scala 416:33]
  wire  _GEN_5758 = invalidate ? _GEN_5242 : _GEN_3694; // @[dcache.scala 416:33]
  wire  _GEN_5759 = invalidate ? _GEN_5243 : _GEN_3695; // @[dcache.scala 416:33]
  wire  _GEN_5760 = invalidate ? _GEN_5244 : _GEN_3696; // @[dcache.scala 416:33]
  wire  _GEN_5761 = invalidate ? _GEN_5245 : _GEN_3697; // @[dcache.scala 416:33]
  wire  _GEN_5762 = invalidate ? _GEN_5246 : _GEN_3698; // @[dcache.scala 416:33]
  wire  _GEN_5763 = invalidate ? _GEN_5247 : _GEN_3699; // @[dcache.scala 416:33]
  wire  _GEN_5764 = invalidate ? _GEN_5248 : _GEN_3700; // @[dcache.scala 416:33]
  wire  _GEN_5765 = invalidate ? _GEN_5249 : _GEN_3701; // @[dcache.scala 416:33]
  wire  _GEN_5766 = invalidate ? _GEN_5250 : _GEN_3702; // @[dcache.scala 416:33]
  wire  _GEN_5767 = invalidate ? _GEN_5251 : _GEN_3703; // @[dcache.scala 416:33]
  wire  _GEN_5768 = invalidate ? _GEN_5252 : _GEN_3704; // @[dcache.scala 416:33]
  wire  _GEN_5769 = invalidate ? _GEN_5253 : _GEN_3705; // @[dcache.scala 416:33]
  wire  _GEN_5770 = invalidate ? _GEN_5254 : _GEN_3706; // @[dcache.scala 416:33]
  wire  _GEN_5771 = invalidate ? _GEN_5255 : _GEN_3707; // @[dcache.scala 416:33]
  wire  _GEN_5772 = invalidate ? _GEN_5256 : _GEN_3708; // @[dcache.scala 416:33]
  wire  _GEN_5773 = invalidate ? _GEN_5257 : _GEN_3709; // @[dcache.scala 416:33]
  wire  _GEN_5774 = invalidate ? _GEN_5258 : _GEN_3710; // @[dcache.scala 416:33]
  wire  _GEN_5775 = invalidate ? _GEN_5259 : _GEN_3711; // @[dcache.scala 416:33]
  wire  _GEN_5776 = invalidate ? _GEN_5260 : _GEN_3712; // @[dcache.scala 416:33]
  wire  _GEN_5777 = invalidate ? _GEN_5261 : _GEN_3713; // @[dcache.scala 416:33]
  wire  _GEN_5778 = invalidate ? _GEN_5262 : _GEN_3714; // @[dcache.scala 416:33]
  wire  _GEN_5779 = invalidate ? _GEN_5263 : _GEN_3715; // @[dcache.scala 416:33]
  wire  _GEN_5780 = invalidate ? _GEN_5264 : _GEN_3716; // @[dcache.scala 416:33]
  wire  _GEN_5781 = invalidate ? _GEN_5265 : _GEN_3717; // @[dcache.scala 416:33]
  wire  _GEN_5782 = invalidate ? _GEN_5266 : _GEN_3718; // @[dcache.scala 416:33]
  wire  _GEN_5783 = invalidate ? _GEN_5267 : _GEN_3719; // @[dcache.scala 416:33]
  wire  _GEN_5784 = invalidate ? _GEN_5268 : _GEN_3720; // @[dcache.scala 416:33]
  wire  _GEN_5785 = invalidate ? _GEN_5269 : _GEN_3721; // @[dcache.scala 416:33]
  wire  _GEN_5786 = invalidate ? _GEN_5270 : _GEN_3722; // @[dcache.scala 416:33]
  wire  _GEN_5787 = invalidate ? _GEN_5271 : _GEN_3723; // @[dcache.scala 416:33]
  wire  _GEN_5788 = invalidate ? _GEN_5272 : _GEN_3724; // @[dcache.scala 416:33]
  wire  _GEN_5789 = invalidate ? _GEN_5273 : _GEN_3725; // @[dcache.scala 416:33]
  wire  _GEN_5790 = invalidate ? _GEN_5274 : _GEN_3726; // @[dcache.scala 416:33]
  wire  _GEN_5791 = invalidate ? _GEN_5275 : _GEN_3727; // @[dcache.scala 416:33]
  wire  _GEN_5792 = invalidate ? _GEN_5276 : _GEN_3728; // @[dcache.scala 416:33]
  wire  _GEN_5793 = invalidate ? _GEN_5277 : _GEN_3729; // @[dcache.scala 416:33]
  wire  _GEN_5794 = invalidate ? _GEN_5278 : _GEN_3730; // @[dcache.scala 416:33]
  wire  _GEN_5795 = invalidate ? _GEN_5279 : _GEN_3731; // @[dcache.scala 416:33]
  wire  _GEN_5796 = invalidate ? _GEN_5280 : _GEN_3732; // @[dcache.scala 416:33]
  wire  _GEN_5797 = invalidate ? _GEN_5281 : _GEN_3733; // @[dcache.scala 416:33]
  wire  _GEN_5798 = invalidate ? _GEN_5282 : _GEN_3734; // @[dcache.scala 416:33]
  wire  _GEN_5799 = invalidate ? _GEN_5283 : _GEN_3735; // @[dcache.scala 416:33]
  wire  _GEN_5800 = invalidate ? _GEN_5284 : _GEN_3736; // @[dcache.scala 416:33]
  wire  _GEN_5801 = invalidate ? _GEN_5285 : _GEN_3737; // @[dcache.scala 416:33]
  wire  _GEN_5802 = invalidate ? _GEN_5286 : _GEN_3738; // @[dcache.scala 416:33]
  wire  _GEN_5803 = invalidate ? _GEN_5287 : _GEN_3739; // @[dcache.scala 416:33]
  wire  _GEN_5804 = invalidate ? _GEN_5288 : _GEN_3740; // @[dcache.scala 416:33]
  wire  _GEN_5805 = invalidate ? _GEN_5289 : _GEN_3741; // @[dcache.scala 416:33]
  wire  _GEN_5806 = invalidate ? _GEN_5290 : _GEN_3742; // @[dcache.scala 416:33]
  wire  _GEN_5807 = invalidate ? _GEN_5291 : _GEN_3743; // @[dcache.scala 416:33]
  wire  _GEN_5808 = invalidate ? _GEN_5292 : _GEN_3744; // @[dcache.scala 416:33]
  wire  _GEN_5809 = invalidate ? _GEN_5293 : _GEN_3745; // @[dcache.scala 416:33]
  wire  _GEN_5810 = invalidate ? _GEN_5294 : _GEN_3746; // @[dcache.scala 416:33]
  wire  _GEN_5811 = invalidate ? _GEN_5295 : _GEN_3747; // @[dcache.scala 416:33]
  wire  _GEN_5812 = invalidate ? _GEN_5296 : _GEN_3748; // @[dcache.scala 416:33]
  wire  _GEN_5813 = invalidate ? _GEN_5297 : _GEN_3749; // @[dcache.scala 416:33]
  wire  _GEN_5814 = invalidate ? _GEN_5298 : _GEN_3750; // @[dcache.scala 416:33]
  wire  _GEN_5815 = invalidate ? _GEN_5299 : _GEN_3751; // @[dcache.scala 416:33]
  wire  _GEN_5816 = invalidate ? _GEN_5300 : _GEN_3752; // @[dcache.scala 416:33]
  wire  _GEN_5817 = invalidate ? _GEN_5301 : _GEN_3753; // @[dcache.scala 416:33]
  wire  _GEN_5818 = invalidate ? _GEN_5302 : _GEN_3754; // @[dcache.scala 416:33]
  wire  _GEN_5819 = invalidate ? _GEN_5303 : _GEN_3755; // @[dcache.scala 416:33]
  wire  _GEN_5820 = invalidate ? _GEN_5304 : _GEN_3756; // @[dcache.scala 416:33]
  wire  _GEN_5821 = invalidate ? _GEN_5305 : _GEN_3757; // @[dcache.scala 416:33]
  wire  _GEN_5822 = invalidate ? _GEN_5306 : _GEN_3758; // @[dcache.scala 416:33]
  wire  _GEN_5823 = invalidate ? _GEN_5307 : _GEN_3759; // @[dcache.scala 416:33]
  wire  _GEN_5824 = invalidate ? _GEN_5308 : _GEN_3760; // @[dcache.scala 416:33]
  wire  _GEN_5825 = invalidate ? _GEN_5309 : _GEN_3761; // @[dcache.scala 416:33]
  wire  _GEN_5826 = invalidate ? _GEN_5310 : _GEN_3762; // @[dcache.scala 416:33]
  wire  _GEN_5827 = invalidate ? _GEN_5311 : _GEN_3763; // @[dcache.scala 416:33]
  wire  _GEN_5828 = invalidate ? _GEN_5312 : _GEN_3764; // @[dcache.scala 416:33]
  wire  _GEN_5829 = invalidate ? _GEN_5313 : _GEN_3765; // @[dcache.scala 416:33]
  wire  _GEN_5830 = invalidate ? _GEN_5314 : _GEN_3766; // @[dcache.scala 416:33]
  wire  _GEN_5831 = invalidate ? _GEN_5315 : _GEN_3767; // @[dcache.scala 416:33]
  wire  _GEN_5832 = invalidate ? _GEN_5316 : _GEN_3768; // @[dcache.scala 416:33]
  wire  _GEN_5833 = invalidate ? _GEN_5317 : _GEN_3769; // @[dcache.scala 416:33]
  wire  _GEN_5834 = invalidate ? _GEN_5318 : _GEN_3770; // @[dcache.scala 416:33]
  wire  _GEN_5835 = invalidate ? _GEN_5319 : _GEN_3771; // @[dcache.scala 416:33]
  wire  _GEN_5836 = invalidate ? _GEN_5320 : _GEN_3772; // @[dcache.scala 416:33]
  wire  _GEN_5837 = invalidate ? _GEN_5321 : _GEN_3773; // @[dcache.scala 416:33]
  wire  _GEN_5838 = invalidate ? _GEN_5322 : _GEN_3774; // @[dcache.scala 416:33]
  wire  _GEN_5839 = invalidate ? _GEN_5323 : _GEN_3775; // @[dcache.scala 416:33]
  wire  _GEN_5840 = invalidate ? _GEN_5324 : _GEN_3776; // @[dcache.scala 416:33]
  wire  _GEN_5841 = invalidate ? _GEN_5325 : _GEN_3777; // @[dcache.scala 416:33]
  wire  _GEN_5842 = invalidate ? _GEN_5326 : _GEN_3778; // @[dcache.scala 416:33]
  wire  _GEN_5843 = invalidate ? _GEN_5327 : _GEN_3779; // @[dcache.scala 416:33]
  wire  _GEN_5844 = invalidate ? _GEN_5328 : _GEN_3780; // @[dcache.scala 416:33]
  wire  _GEN_5845 = invalidate ? _GEN_5329 : _GEN_3781; // @[dcache.scala 416:33]
  wire  _GEN_5846 = invalidate ? _GEN_5330 : _GEN_3782; // @[dcache.scala 416:33]
  wire  _GEN_5847 = invalidate ? _GEN_5331 : _GEN_3783; // @[dcache.scala 416:33]
  wire  _GEN_5848 = invalidate ? _GEN_5332 : _GEN_3784; // @[dcache.scala 416:33]
  wire  _GEN_5849 = invalidate ? _GEN_5333 : _GEN_3785; // @[dcache.scala 416:33]
  wire  _GEN_5850 = invalidate ? _GEN_5334 : _GEN_3786; // @[dcache.scala 416:33]
  wire  _GEN_5851 = invalidate ? _GEN_5335 : _GEN_3787; // @[dcache.scala 416:33]
  wire  _GEN_5852 = invalidate ? _GEN_5336 : _GEN_3788; // @[dcache.scala 416:33]
  wire  _GEN_5853 = invalidate ? _GEN_5337 : _GEN_3789; // @[dcache.scala 416:33]
  wire  _GEN_5854 = invalidate ? _GEN_5338 : _GEN_3790; // @[dcache.scala 416:33]
  wire  _GEN_5855 = invalidate ? _GEN_5339 : _GEN_3791; // @[dcache.scala 416:33]
  wire  _GEN_5856 = invalidate ? _GEN_5340 : _GEN_3792; // @[dcache.scala 416:33]
  wire  _GEN_5857 = invalidate ? _GEN_5341 : _GEN_3793; // @[dcache.scala 416:33]
  wire  _GEN_5858 = invalidate ? _GEN_5342 : _GEN_3794; // @[dcache.scala 416:33]
  wire  _GEN_5859 = invalidate ? _GEN_5343 : _GEN_3795; // @[dcache.scala 416:33]
  wire  _GEN_5860 = invalidate ? _GEN_5344 : _GEN_3796; // @[dcache.scala 416:33]
  wire  _GEN_5861 = invalidate ? _GEN_5345 : _GEN_3797; // @[dcache.scala 416:33]
  wire  _GEN_5862 = invalidate ? _GEN_5346 : _GEN_3798; // @[dcache.scala 416:33]
  wire  _GEN_5863 = invalidate ? _GEN_5347 : _GEN_3799; // @[dcache.scala 416:33]
  wire  _GEN_5864 = invalidate ? _GEN_5348 : _GEN_3800; // @[dcache.scala 416:33]
  wire  _GEN_5865 = invalidate ? _GEN_5349 : _GEN_3801; // @[dcache.scala 416:33]
  wire  _GEN_5866 = invalidate ? _GEN_5350 : _GEN_3802; // @[dcache.scala 416:33]
  wire  _GEN_5867 = invalidate ? _GEN_5351 : _GEN_3803; // @[dcache.scala 416:33]
  wire  _GEN_5868 = invalidate ? _GEN_5352 : _GEN_3804; // @[dcache.scala 416:33]
  wire  _GEN_5869 = invalidate ? _GEN_5353 : _GEN_3805; // @[dcache.scala 416:33]
  wire  _GEN_5870 = invalidate ? _GEN_5354 : _GEN_3806; // @[dcache.scala 416:33]
  wire  _GEN_5871 = invalidate ? _GEN_5355 : _GEN_3807; // @[dcache.scala 416:33]
  wire  _GEN_5872 = invalidate ? _GEN_5356 : _GEN_3808; // @[dcache.scala 416:33]
  wire  _GEN_5873 = invalidate ? _GEN_5357 : _GEN_3809; // @[dcache.scala 416:33]
  wire  _GEN_5874 = invalidate ? _GEN_5358 : _GEN_3810; // @[dcache.scala 416:33]
  wire  _GEN_5875 = invalidate ? _GEN_5359 : _GEN_3811; // @[dcache.scala 416:33]
  wire  _GEN_5876 = invalidate ? _GEN_5360 : _GEN_3812; // @[dcache.scala 416:33]
  wire  _GEN_5877 = invalidate ? _GEN_5361 : _GEN_3813; // @[dcache.scala 416:33]
  wire  _GEN_5878 = invalidate ? _GEN_5362 : _GEN_3814; // @[dcache.scala 416:33]
  wire  _GEN_5879 = invalidate ? _GEN_5363 : _GEN_3815; // @[dcache.scala 416:33]
  wire  _GEN_5880 = invalidate ? _GEN_5364 : _GEN_3816; // @[dcache.scala 416:33]
  wire  _GEN_5881 = invalidate ? _GEN_5365 : _GEN_3817; // @[dcache.scala 416:33]
  wire  _GEN_5882 = invalidate ? _GEN_5366 : _GEN_3818; // @[dcache.scala 416:33]
  wire  _GEN_5883 = invalidate ? _GEN_5367 : _GEN_3819; // @[dcache.scala 416:33]
  wire  _GEN_5884 = invalidate ? _GEN_5368 : _GEN_3820; // @[dcache.scala 416:33]
  wire  _GEN_5885 = invalidate ? _GEN_5369 : _GEN_3821; // @[dcache.scala 416:33]
  wire  _GEN_5886 = invalidate ? _GEN_5370 : _GEN_3822; // @[dcache.scala 416:33]
  wire  _GEN_5887 = invalidate ? _GEN_5371 : _GEN_3823; // @[dcache.scala 416:33]
  wire  _GEN_5888 = invalidate ? _GEN_5372 : _GEN_3824; // @[dcache.scala 416:33]
  wire  _GEN_5889 = invalidate ? _GEN_5373 : _GEN_3825; // @[dcache.scala 416:33]
  wire  _GEN_5890 = invalidate ? _GEN_5374 : _GEN_3826; // @[dcache.scala 416:33]
  wire  _GEN_5891 = invalidate ? _GEN_5375 : _GEN_3827; // @[dcache.scala 416:33]
  wire  _GEN_5892 = invalidate ? _GEN_5376 : _GEN_3828; // @[dcache.scala 416:33]
  wire  _GEN_5893 = invalidate ? _GEN_5377 : _GEN_3829; // @[dcache.scala 416:33]
  wire  _GEN_5894 = invalidate ? _GEN_5378 : _GEN_3830; // @[dcache.scala 416:33]
  wire  _GEN_5895 = invalidate ? _GEN_5379 : _GEN_3831; // @[dcache.scala 416:33]
  wire  _GEN_5896 = invalidate ? _GEN_5380 : _GEN_3832; // @[dcache.scala 416:33]
  wire  _GEN_5897 = invalidate ? _GEN_5381 : _GEN_3833; // @[dcache.scala 416:33]
  wire  _GEN_5898 = invalidate ? _GEN_5382 : _GEN_3834; // @[dcache.scala 416:33]
  wire  _GEN_5899 = invalidate ? _GEN_5383 : _GEN_3835; // @[dcache.scala 416:33]
  wire  _GEN_5900 = invalidate ? _GEN_5384 : _GEN_3836; // @[dcache.scala 416:33]
  wire  _GEN_5901 = invalidate ? _GEN_5385 : _GEN_3837; // @[dcache.scala 416:33]
  wire  _GEN_5902 = invalidate ? _GEN_5386 : _GEN_3838; // @[dcache.scala 416:33]
  wire  _GEN_5903 = invalidate ? _GEN_5387 : _GEN_3839; // @[dcache.scala 416:33]
  wire  _GEN_5904 = invalidate ? _GEN_5388 : _GEN_3840; // @[dcache.scala 416:33]
  wire  _GEN_5905 = invalidate ? _GEN_5389 : _GEN_3841; // @[dcache.scala 416:33]
  wire  _GEN_5906 = invalidate ? _GEN_5390 : _GEN_3842; // @[dcache.scala 416:33]
  wire  _GEN_5907 = invalidate ? _GEN_5391 : _GEN_3843; // @[dcache.scala 416:33]
  wire  _GEN_5908 = invalidate ? _GEN_5392 : _GEN_3844; // @[dcache.scala 416:33]
  wire  _GEN_5909 = invalidate ? _GEN_5393 : _GEN_3845; // @[dcache.scala 416:33]
  wire  _GEN_5910 = invalidate ? _GEN_5394 : _GEN_3846; // @[dcache.scala 416:33]
  wire  _GEN_5911 = invalidate ? _GEN_5395 : _GEN_3847; // @[dcache.scala 416:33]
  wire  _GEN_5912 = invalidate ? _GEN_5396 : _GEN_3848; // @[dcache.scala 416:33]
  wire  _GEN_5913 = invalidate ? _GEN_5397 : _GEN_3849; // @[dcache.scala 416:33]
  wire  _GEN_5914 = invalidate ? _GEN_5398 : _GEN_3850; // @[dcache.scala 416:33]
  wire  _GEN_5915 = _T_7 & _T_51; // @[dcache.scala 157:25 397:36]
  wire [31:0] _GEN_5916 = _T_7 ? _GEN_2301 : 32'h7777; // @[dcache.scala 155:25 397:36]
  wire [2:0] _GEN_5917 = _T_7 ? _GEN_2302 : 3'h0; // @[dcache.scala 397:36 406:61]
  wire  _GEN_5918 = _T_7 ? _GEN_2303 : req_valid; // @[dcache.scala 116:34 397:36]
  wire  _GEN_5919 = _T_7 ? 1'h0 : 1'h1; // @[dcache.scala 397:36 97:21 407:61]
  wire [21:0] _GEN_5920 = _T_7 ? 22'h0 : _GEN_2818; // @[dcache.scala 397:36 98:21]
  wire [20:0] _GEN_5921 = _T_7 ? 21'h0 : _GEN_5399; // @[dcache.scala 143:25 397:36]
  wire [20:0] _GEN_5922 = _T_7 ? 21'h0 : _GEN_5400; // @[dcache.scala 143:25 397:36]
  wire  _GEN_5923 = _T_7 ? 1'h0 : _GEN_5401; // @[dcache.scala 144:25 397:36]
  wire  _GEN_5924 = _T_7 ? 1'h0 : _GEN_5402; // @[dcache.scala 144:25 397:36]
  wire  _GEN_5925 = _T_7 ? dirty_0_0 : _GEN_5403; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5926 = _T_7 ? dirty_0_1 : _GEN_5404; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5927 = _T_7 ? dirty_0_2 : _GEN_5405; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5928 = _T_7 ? dirty_0_3 : _GEN_5406; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5929 = _T_7 ? dirty_0_4 : _GEN_5407; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5930 = _T_7 ? dirty_0_5 : _GEN_5408; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5931 = _T_7 ? dirty_0_6 : _GEN_5409; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5932 = _T_7 ? dirty_0_7 : _GEN_5410; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5933 = _T_7 ? dirty_0_8 : _GEN_5411; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5934 = _T_7 ? dirty_0_9 : _GEN_5412; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5935 = _T_7 ? dirty_0_10 : _GEN_5413; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5936 = _T_7 ? dirty_0_11 : _GEN_5414; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5937 = _T_7 ? dirty_0_12 : _GEN_5415; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5938 = _T_7 ? dirty_0_13 : _GEN_5416; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5939 = _T_7 ? dirty_0_14 : _GEN_5417; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5940 = _T_7 ? dirty_0_15 : _GEN_5418; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5941 = _T_7 ? dirty_0_16 : _GEN_5419; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5942 = _T_7 ? dirty_0_17 : _GEN_5420; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5943 = _T_7 ? dirty_0_18 : _GEN_5421; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5944 = _T_7 ? dirty_0_19 : _GEN_5422; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5945 = _T_7 ? dirty_0_20 : _GEN_5423; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5946 = _T_7 ? dirty_0_21 : _GEN_5424; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5947 = _T_7 ? dirty_0_22 : _GEN_5425; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5948 = _T_7 ? dirty_0_23 : _GEN_5426; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5949 = _T_7 ? dirty_0_24 : _GEN_5427; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5950 = _T_7 ? dirty_0_25 : _GEN_5428; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5951 = _T_7 ? dirty_0_26 : _GEN_5429; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5952 = _T_7 ? dirty_0_27 : _GEN_5430; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5953 = _T_7 ? dirty_0_28 : _GEN_5431; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5954 = _T_7 ? dirty_0_29 : _GEN_5432; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5955 = _T_7 ? dirty_0_30 : _GEN_5433; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5956 = _T_7 ? dirty_0_31 : _GEN_5434; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5957 = _T_7 ? dirty_0_32 : _GEN_5435; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5958 = _T_7 ? dirty_0_33 : _GEN_5436; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5959 = _T_7 ? dirty_0_34 : _GEN_5437; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5960 = _T_7 ? dirty_0_35 : _GEN_5438; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5961 = _T_7 ? dirty_0_36 : _GEN_5439; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5962 = _T_7 ? dirty_0_37 : _GEN_5440; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5963 = _T_7 ? dirty_0_38 : _GEN_5441; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5964 = _T_7 ? dirty_0_39 : _GEN_5442; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5965 = _T_7 ? dirty_0_40 : _GEN_5443; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5966 = _T_7 ? dirty_0_41 : _GEN_5444; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5967 = _T_7 ? dirty_0_42 : _GEN_5445; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5968 = _T_7 ? dirty_0_43 : _GEN_5446; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5969 = _T_7 ? dirty_0_44 : _GEN_5447; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5970 = _T_7 ? dirty_0_45 : _GEN_5448; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5971 = _T_7 ? dirty_0_46 : _GEN_5449; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5972 = _T_7 ? dirty_0_47 : _GEN_5450; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5973 = _T_7 ? dirty_0_48 : _GEN_5451; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5974 = _T_7 ? dirty_0_49 : _GEN_5452; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5975 = _T_7 ? dirty_0_50 : _GEN_5453; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5976 = _T_7 ? dirty_0_51 : _GEN_5454; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5977 = _T_7 ? dirty_0_52 : _GEN_5455; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5978 = _T_7 ? dirty_0_53 : _GEN_5456; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5979 = _T_7 ? dirty_0_54 : _GEN_5457; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5980 = _T_7 ? dirty_0_55 : _GEN_5458; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5981 = _T_7 ? dirty_0_56 : _GEN_5459; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5982 = _T_7 ? dirty_0_57 : _GEN_5460; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5983 = _T_7 ? dirty_0_58 : _GEN_5461; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5984 = _T_7 ? dirty_0_59 : _GEN_5462; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5985 = _T_7 ? dirty_0_60 : _GEN_5463; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5986 = _T_7 ? dirty_0_61 : _GEN_5464; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5987 = _T_7 ? dirty_0_62 : _GEN_5465; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5988 = _T_7 ? dirty_0_63 : _GEN_5466; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5989 = _T_7 ? dirty_0_64 : _GEN_5467; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5990 = _T_7 ? dirty_0_65 : _GEN_5468; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5991 = _T_7 ? dirty_0_66 : _GEN_5469; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5992 = _T_7 ? dirty_0_67 : _GEN_5470; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5993 = _T_7 ? dirty_0_68 : _GEN_5471; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5994 = _T_7 ? dirty_0_69 : _GEN_5472; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5995 = _T_7 ? dirty_0_70 : _GEN_5473; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5996 = _T_7 ? dirty_0_71 : _GEN_5474; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5997 = _T_7 ? dirty_0_72 : _GEN_5475; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5998 = _T_7 ? dirty_0_73 : _GEN_5476; // @[dcache.scala 113:28 397:36]
  wire  _GEN_5999 = _T_7 ? dirty_0_74 : _GEN_5477; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6000 = _T_7 ? dirty_0_75 : _GEN_5478; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6001 = _T_7 ? dirty_0_76 : _GEN_5479; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6002 = _T_7 ? dirty_0_77 : _GEN_5480; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6003 = _T_7 ? dirty_0_78 : _GEN_5481; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6004 = _T_7 ? dirty_0_79 : _GEN_5482; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6005 = _T_7 ? dirty_0_80 : _GEN_5483; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6006 = _T_7 ? dirty_0_81 : _GEN_5484; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6007 = _T_7 ? dirty_0_82 : _GEN_5485; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6008 = _T_7 ? dirty_0_83 : _GEN_5486; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6009 = _T_7 ? dirty_0_84 : _GEN_5487; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6010 = _T_7 ? dirty_0_85 : _GEN_5488; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6011 = _T_7 ? dirty_0_86 : _GEN_5489; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6012 = _T_7 ? dirty_0_87 : _GEN_5490; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6013 = _T_7 ? dirty_0_88 : _GEN_5491; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6014 = _T_7 ? dirty_0_89 : _GEN_5492; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6015 = _T_7 ? dirty_0_90 : _GEN_5493; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6016 = _T_7 ? dirty_0_91 : _GEN_5494; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6017 = _T_7 ? dirty_0_92 : _GEN_5495; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6018 = _T_7 ? dirty_0_93 : _GEN_5496; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6019 = _T_7 ? dirty_0_94 : _GEN_5497; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6020 = _T_7 ? dirty_0_95 : _GEN_5498; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6021 = _T_7 ? dirty_0_96 : _GEN_5499; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6022 = _T_7 ? dirty_0_97 : _GEN_5500; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6023 = _T_7 ? dirty_0_98 : _GEN_5501; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6024 = _T_7 ? dirty_0_99 : _GEN_5502; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6025 = _T_7 ? dirty_0_100 : _GEN_5503; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6026 = _T_7 ? dirty_0_101 : _GEN_5504; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6027 = _T_7 ? dirty_0_102 : _GEN_5505; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6028 = _T_7 ? dirty_0_103 : _GEN_5506; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6029 = _T_7 ? dirty_0_104 : _GEN_5507; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6030 = _T_7 ? dirty_0_105 : _GEN_5508; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6031 = _T_7 ? dirty_0_106 : _GEN_5509; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6032 = _T_7 ? dirty_0_107 : _GEN_5510; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6033 = _T_7 ? dirty_0_108 : _GEN_5511; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6034 = _T_7 ? dirty_0_109 : _GEN_5512; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6035 = _T_7 ? dirty_0_110 : _GEN_5513; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6036 = _T_7 ? dirty_0_111 : _GEN_5514; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6037 = _T_7 ? dirty_0_112 : _GEN_5515; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6038 = _T_7 ? dirty_0_113 : _GEN_5516; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6039 = _T_7 ? dirty_0_114 : _GEN_5517; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6040 = _T_7 ? dirty_0_115 : _GEN_5518; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6041 = _T_7 ? dirty_0_116 : _GEN_5519; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6042 = _T_7 ? dirty_0_117 : _GEN_5520; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6043 = _T_7 ? dirty_0_118 : _GEN_5521; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6044 = _T_7 ? dirty_0_119 : _GEN_5522; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6045 = _T_7 ? dirty_0_120 : _GEN_5523; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6046 = _T_7 ? dirty_0_121 : _GEN_5524; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6047 = _T_7 ? dirty_0_122 : _GEN_5525; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6048 = _T_7 ? dirty_0_123 : _GEN_5526; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6049 = _T_7 ? dirty_0_124 : _GEN_5527; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6050 = _T_7 ? dirty_0_125 : _GEN_5528; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6051 = _T_7 ? dirty_0_126 : _GEN_5529; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6052 = _T_7 ? dirty_0_127 : _GEN_5530; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6053 = _T_7 ? dirty_0_128 : _GEN_5531; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6054 = _T_7 ? dirty_0_129 : _GEN_5532; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6055 = _T_7 ? dirty_0_130 : _GEN_5533; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6056 = _T_7 ? dirty_0_131 : _GEN_5534; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6057 = _T_7 ? dirty_0_132 : _GEN_5535; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6058 = _T_7 ? dirty_0_133 : _GEN_5536; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6059 = _T_7 ? dirty_0_134 : _GEN_5537; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6060 = _T_7 ? dirty_0_135 : _GEN_5538; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6061 = _T_7 ? dirty_0_136 : _GEN_5539; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6062 = _T_7 ? dirty_0_137 : _GEN_5540; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6063 = _T_7 ? dirty_0_138 : _GEN_5541; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6064 = _T_7 ? dirty_0_139 : _GEN_5542; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6065 = _T_7 ? dirty_0_140 : _GEN_5543; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6066 = _T_7 ? dirty_0_141 : _GEN_5544; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6067 = _T_7 ? dirty_0_142 : _GEN_5545; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6068 = _T_7 ? dirty_0_143 : _GEN_5546; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6069 = _T_7 ? dirty_0_144 : _GEN_5547; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6070 = _T_7 ? dirty_0_145 : _GEN_5548; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6071 = _T_7 ? dirty_0_146 : _GEN_5549; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6072 = _T_7 ? dirty_0_147 : _GEN_5550; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6073 = _T_7 ? dirty_0_148 : _GEN_5551; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6074 = _T_7 ? dirty_0_149 : _GEN_5552; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6075 = _T_7 ? dirty_0_150 : _GEN_5553; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6076 = _T_7 ? dirty_0_151 : _GEN_5554; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6077 = _T_7 ? dirty_0_152 : _GEN_5555; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6078 = _T_7 ? dirty_0_153 : _GEN_5556; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6079 = _T_7 ? dirty_0_154 : _GEN_5557; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6080 = _T_7 ? dirty_0_155 : _GEN_5558; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6081 = _T_7 ? dirty_0_156 : _GEN_5559; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6082 = _T_7 ? dirty_0_157 : _GEN_5560; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6083 = _T_7 ? dirty_0_158 : _GEN_5561; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6084 = _T_7 ? dirty_0_159 : _GEN_5562; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6085 = _T_7 ? dirty_0_160 : _GEN_5563; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6086 = _T_7 ? dirty_0_161 : _GEN_5564; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6087 = _T_7 ? dirty_0_162 : _GEN_5565; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6088 = _T_7 ? dirty_0_163 : _GEN_5566; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6089 = _T_7 ? dirty_0_164 : _GEN_5567; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6090 = _T_7 ? dirty_0_165 : _GEN_5568; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6091 = _T_7 ? dirty_0_166 : _GEN_5569; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6092 = _T_7 ? dirty_0_167 : _GEN_5570; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6093 = _T_7 ? dirty_0_168 : _GEN_5571; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6094 = _T_7 ? dirty_0_169 : _GEN_5572; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6095 = _T_7 ? dirty_0_170 : _GEN_5573; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6096 = _T_7 ? dirty_0_171 : _GEN_5574; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6097 = _T_7 ? dirty_0_172 : _GEN_5575; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6098 = _T_7 ? dirty_0_173 : _GEN_5576; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6099 = _T_7 ? dirty_0_174 : _GEN_5577; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6100 = _T_7 ? dirty_0_175 : _GEN_5578; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6101 = _T_7 ? dirty_0_176 : _GEN_5579; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6102 = _T_7 ? dirty_0_177 : _GEN_5580; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6103 = _T_7 ? dirty_0_178 : _GEN_5581; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6104 = _T_7 ? dirty_0_179 : _GEN_5582; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6105 = _T_7 ? dirty_0_180 : _GEN_5583; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6106 = _T_7 ? dirty_0_181 : _GEN_5584; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6107 = _T_7 ? dirty_0_182 : _GEN_5585; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6108 = _T_7 ? dirty_0_183 : _GEN_5586; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6109 = _T_7 ? dirty_0_184 : _GEN_5587; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6110 = _T_7 ? dirty_0_185 : _GEN_5588; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6111 = _T_7 ? dirty_0_186 : _GEN_5589; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6112 = _T_7 ? dirty_0_187 : _GEN_5590; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6113 = _T_7 ? dirty_0_188 : _GEN_5591; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6114 = _T_7 ? dirty_0_189 : _GEN_5592; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6115 = _T_7 ? dirty_0_190 : _GEN_5593; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6116 = _T_7 ? dirty_0_191 : _GEN_5594; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6117 = _T_7 ? dirty_0_192 : _GEN_5595; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6118 = _T_7 ? dirty_0_193 : _GEN_5596; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6119 = _T_7 ? dirty_0_194 : _GEN_5597; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6120 = _T_7 ? dirty_0_195 : _GEN_5598; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6121 = _T_7 ? dirty_0_196 : _GEN_5599; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6122 = _T_7 ? dirty_0_197 : _GEN_5600; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6123 = _T_7 ? dirty_0_198 : _GEN_5601; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6124 = _T_7 ? dirty_0_199 : _GEN_5602; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6125 = _T_7 ? dirty_0_200 : _GEN_5603; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6126 = _T_7 ? dirty_0_201 : _GEN_5604; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6127 = _T_7 ? dirty_0_202 : _GEN_5605; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6128 = _T_7 ? dirty_0_203 : _GEN_5606; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6129 = _T_7 ? dirty_0_204 : _GEN_5607; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6130 = _T_7 ? dirty_0_205 : _GEN_5608; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6131 = _T_7 ? dirty_0_206 : _GEN_5609; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6132 = _T_7 ? dirty_0_207 : _GEN_5610; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6133 = _T_7 ? dirty_0_208 : _GEN_5611; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6134 = _T_7 ? dirty_0_209 : _GEN_5612; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6135 = _T_7 ? dirty_0_210 : _GEN_5613; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6136 = _T_7 ? dirty_0_211 : _GEN_5614; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6137 = _T_7 ? dirty_0_212 : _GEN_5615; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6138 = _T_7 ? dirty_0_213 : _GEN_5616; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6139 = _T_7 ? dirty_0_214 : _GEN_5617; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6140 = _T_7 ? dirty_0_215 : _GEN_5618; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6141 = _T_7 ? dirty_0_216 : _GEN_5619; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6142 = _T_7 ? dirty_0_217 : _GEN_5620; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6143 = _T_7 ? dirty_0_218 : _GEN_5621; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6144 = _T_7 ? dirty_0_219 : _GEN_5622; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6145 = _T_7 ? dirty_0_220 : _GEN_5623; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6146 = _T_7 ? dirty_0_221 : _GEN_5624; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6147 = _T_7 ? dirty_0_222 : _GEN_5625; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6148 = _T_7 ? dirty_0_223 : _GEN_5626; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6149 = _T_7 ? dirty_0_224 : _GEN_5627; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6150 = _T_7 ? dirty_0_225 : _GEN_5628; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6151 = _T_7 ? dirty_0_226 : _GEN_5629; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6152 = _T_7 ? dirty_0_227 : _GEN_5630; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6153 = _T_7 ? dirty_0_228 : _GEN_5631; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6154 = _T_7 ? dirty_0_229 : _GEN_5632; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6155 = _T_7 ? dirty_0_230 : _GEN_5633; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6156 = _T_7 ? dirty_0_231 : _GEN_5634; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6157 = _T_7 ? dirty_0_232 : _GEN_5635; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6158 = _T_7 ? dirty_0_233 : _GEN_5636; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6159 = _T_7 ? dirty_0_234 : _GEN_5637; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6160 = _T_7 ? dirty_0_235 : _GEN_5638; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6161 = _T_7 ? dirty_0_236 : _GEN_5639; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6162 = _T_7 ? dirty_0_237 : _GEN_5640; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6163 = _T_7 ? dirty_0_238 : _GEN_5641; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6164 = _T_7 ? dirty_0_239 : _GEN_5642; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6165 = _T_7 ? dirty_0_240 : _GEN_5643; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6166 = _T_7 ? dirty_0_241 : _GEN_5644; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6167 = _T_7 ? dirty_0_242 : _GEN_5645; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6168 = _T_7 ? dirty_0_243 : _GEN_5646; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6169 = _T_7 ? dirty_0_244 : _GEN_5647; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6170 = _T_7 ? dirty_0_245 : _GEN_5648; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6171 = _T_7 ? dirty_0_246 : _GEN_5649; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6172 = _T_7 ? dirty_0_247 : _GEN_5650; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6173 = _T_7 ? dirty_0_248 : _GEN_5651; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6174 = _T_7 ? dirty_0_249 : _GEN_5652; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6175 = _T_7 ? dirty_0_250 : _GEN_5653; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6176 = _T_7 ? dirty_0_251 : _GEN_5654; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6177 = _T_7 ? dirty_0_252 : _GEN_5655; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6178 = _T_7 ? dirty_0_253 : _GEN_5656; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6179 = _T_7 ? dirty_0_254 : _GEN_5657; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6180 = _T_7 ? dirty_0_255 : _GEN_5658; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6181 = _T_7 ? dirty_1_0 : _GEN_5659; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6182 = _T_7 ? dirty_1_1 : _GEN_5660; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6183 = _T_7 ? dirty_1_2 : _GEN_5661; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6184 = _T_7 ? dirty_1_3 : _GEN_5662; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6185 = _T_7 ? dirty_1_4 : _GEN_5663; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6186 = _T_7 ? dirty_1_5 : _GEN_5664; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6187 = _T_7 ? dirty_1_6 : _GEN_5665; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6188 = _T_7 ? dirty_1_7 : _GEN_5666; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6189 = _T_7 ? dirty_1_8 : _GEN_5667; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6190 = _T_7 ? dirty_1_9 : _GEN_5668; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6191 = _T_7 ? dirty_1_10 : _GEN_5669; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6192 = _T_7 ? dirty_1_11 : _GEN_5670; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6193 = _T_7 ? dirty_1_12 : _GEN_5671; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6194 = _T_7 ? dirty_1_13 : _GEN_5672; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6195 = _T_7 ? dirty_1_14 : _GEN_5673; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6196 = _T_7 ? dirty_1_15 : _GEN_5674; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6197 = _T_7 ? dirty_1_16 : _GEN_5675; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6198 = _T_7 ? dirty_1_17 : _GEN_5676; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6199 = _T_7 ? dirty_1_18 : _GEN_5677; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6200 = _T_7 ? dirty_1_19 : _GEN_5678; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6201 = _T_7 ? dirty_1_20 : _GEN_5679; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6202 = _T_7 ? dirty_1_21 : _GEN_5680; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6203 = _T_7 ? dirty_1_22 : _GEN_5681; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6204 = _T_7 ? dirty_1_23 : _GEN_5682; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6205 = _T_7 ? dirty_1_24 : _GEN_5683; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6206 = _T_7 ? dirty_1_25 : _GEN_5684; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6207 = _T_7 ? dirty_1_26 : _GEN_5685; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6208 = _T_7 ? dirty_1_27 : _GEN_5686; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6209 = _T_7 ? dirty_1_28 : _GEN_5687; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6210 = _T_7 ? dirty_1_29 : _GEN_5688; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6211 = _T_7 ? dirty_1_30 : _GEN_5689; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6212 = _T_7 ? dirty_1_31 : _GEN_5690; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6213 = _T_7 ? dirty_1_32 : _GEN_5691; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6214 = _T_7 ? dirty_1_33 : _GEN_5692; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6215 = _T_7 ? dirty_1_34 : _GEN_5693; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6216 = _T_7 ? dirty_1_35 : _GEN_5694; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6217 = _T_7 ? dirty_1_36 : _GEN_5695; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6218 = _T_7 ? dirty_1_37 : _GEN_5696; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6219 = _T_7 ? dirty_1_38 : _GEN_5697; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6220 = _T_7 ? dirty_1_39 : _GEN_5698; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6221 = _T_7 ? dirty_1_40 : _GEN_5699; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6222 = _T_7 ? dirty_1_41 : _GEN_5700; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6223 = _T_7 ? dirty_1_42 : _GEN_5701; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6224 = _T_7 ? dirty_1_43 : _GEN_5702; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6225 = _T_7 ? dirty_1_44 : _GEN_5703; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6226 = _T_7 ? dirty_1_45 : _GEN_5704; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6227 = _T_7 ? dirty_1_46 : _GEN_5705; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6228 = _T_7 ? dirty_1_47 : _GEN_5706; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6229 = _T_7 ? dirty_1_48 : _GEN_5707; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6230 = _T_7 ? dirty_1_49 : _GEN_5708; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6231 = _T_7 ? dirty_1_50 : _GEN_5709; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6232 = _T_7 ? dirty_1_51 : _GEN_5710; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6233 = _T_7 ? dirty_1_52 : _GEN_5711; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6234 = _T_7 ? dirty_1_53 : _GEN_5712; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6235 = _T_7 ? dirty_1_54 : _GEN_5713; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6236 = _T_7 ? dirty_1_55 : _GEN_5714; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6237 = _T_7 ? dirty_1_56 : _GEN_5715; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6238 = _T_7 ? dirty_1_57 : _GEN_5716; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6239 = _T_7 ? dirty_1_58 : _GEN_5717; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6240 = _T_7 ? dirty_1_59 : _GEN_5718; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6241 = _T_7 ? dirty_1_60 : _GEN_5719; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6242 = _T_7 ? dirty_1_61 : _GEN_5720; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6243 = _T_7 ? dirty_1_62 : _GEN_5721; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6244 = _T_7 ? dirty_1_63 : _GEN_5722; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6245 = _T_7 ? dirty_1_64 : _GEN_5723; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6246 = _T_7 ? dirty_1_65 : _GEN_5724; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6247 = _T_7 ? dirty_1_66 : _GEN_5725; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6248 = _T_7 ? dirty_1_67 : _GEN_5726; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6249 = _T_7 ? dirty_1_68 : _GEN_5727; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6250 = _T_7 ? dirty_1_69 : _GEN_5728; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6251 = _T_7 ? dirty_1_70 : _GEN_5729; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6252 = _T_7 ? dirty_1_71 : _GEN_5730; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6253 = _T_7 ? dirty_1_72 : _GEN_5731; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6254 = _T_7 ? dirty_1_73 : _GEN_5732; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6255 = _T_7 ? dirty_1_74 : _GEN_5733; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6256 = _T_7 ? dirty_1_75 : _GEN_5734; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6257 = _T_7 ? dirty_1_76 : _GEN_5735; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6258 = _T_7 ? dirty_1_77 : _GEN_5736; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6259 = _T_7 ? dirty_1_78 : _GEN_5737; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6260 = _T_7 ? dirty_1_79 : _GEN_5738; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6261 = _T_7 ? dirty_1_80 : _GEN_5739; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6262 = _T_7 ? dirty_1_81 : _GEN_5740; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6263 = _T_7 ? dirty_1_82 : _GEN_5741; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6264 = _T_7 ? dirty_1_83 : _GEN_5742; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6265 = _T_7 ? dirty_1_84 : _GEN_5743; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6266 = _T_7 ? dirty_1_85 : _GEN_5744; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6267 = _T_7 ? dirty_1_86 : _GEN_5745; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6268 = _T_7 ? dirty_1_87 : _GEN_5746; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6269 = _T_7 ? dirty_1_88 : _GEN_5747; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6270 = _T_7 ? dirty_1_89 : _GEN_5748; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6271 = _T_7 ? dirty_1_90 : _GEN_5749; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6272 = _T_7 ? dirty_1_91 : _GEN_5750; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6273 = _T_7 ? dirty_1_92 : _GEN_5751; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6274 = _T_7 ? dirty_1_93 : _GEN_5752; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6275 = _T_7 ? dirty_1_94 : _GEN_5753; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6276 = _T_7 ? dirty_1_95 : _GEN_5754; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6277 = _T_7 ? dirty_1_96 : _GEN_5755; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6278 = _T_7 ? dirty_1_97 : _GEN_5756; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6279 = _T_7 ? dirty_1_98 : _GEN_5757; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6280 = _T_7 ? dirty_1_99 : _GEN_5758; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6281 = _T_7 ? dirty_1_100 : _GEN_5759; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6282 = _T_7 ? dirty_1_101 : _GEN_5760; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6283 = _T_7 ? dirty_1_102 : _GEN_5761; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6284 = _T_7 ? dirty_1_103 : _GEN_5762; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6285 = _T_7 ? dirty_1_104 : _GEN_5763; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6286 = _T_7 ? dirty_1_105 : _GEN_5764; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6287 = _T_7 ? dirty_1_106 : _GEN_5765; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6288 = _T_7 ? dirty_1_107 : _GEN_5766; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6289 = _T_7 ? dirty_1_108 : _GEN_5767; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6290 = _T_7 ? dirty_1_109 : _GEN_5768; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6291 = _T_7 ? dirty_1_110 : _GEN_5769; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6292 = _T_7 ? dirty_1_111 : _GEN_5770; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6293 = _T_7 ? dirty_1_112 : _GEN_5771; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6294 = _T_7 ? dirty_1_113 : _GEN_5772; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6295 = _T_7 ? dirty_1_114 : _GEN_5773; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6296 = _T_7 ? dirty_1_115 : _GEN_5774; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6297 = _T_7 ? dirty_1_116 : _GEN_5775; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6298 = _T_7 ? dirty_1_117 : _GEN_5776; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6299 = _T_7 ? dirty_1_118 : _GEN_5777; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6300 = _T_7 ? dirty_1_119 : _GEN_5778; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6301 = _T_7 ? dirty_1_120 : _GEN_5779; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6302 = _T_7 ? dirty_1_121 : _GEN_5780; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6303 = _T_7 ? dirty_1_122 : _GEN_5781; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6304 = _T_7 ? dirty_1_123 : _GEN_5782; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6305 = _T_7 ? dirty_1_124 : _GEN_5783; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6306 = _T_7 ? dirty_1_125 : _GEN_5784; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6307 = _T_7 ? dirty_1_126 : _GEN_5785; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6308 = _T_7 ? dirty_1_127 : _GEN_5786; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6309 = _T_7 ? dirty_1_128 : _GEN_5787; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6310 = _T_7 ? dirty_1_129 : _GEN_5788; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6311 = _T_7 ? dirty_1_130 : _GEN_5789; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6312 = _T_7 ? dirty_1_131 : _GEN_5790; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6313 = _T_7 ? dirty_1_132 : _GEN_5791; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6314 = _T_7 ? dirty_1_133 : _GEN_5792; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6315 = _T_7 ? dirty_1_134 : _GEN_5793; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6316 = _T_7 ? dirty_1_135 : _GEN_5794; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6317 = _T_7 ? dirty_1_136 : _GEN_5795; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6318 = _T_7 ? dirty_1_137 : _GEN_5796; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6319 = _T_7 ? dirty_1_138 : _GEN_5797; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6320 = _T_7 ? dirty_1_139 : _GEN_5798; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6321 = _T_7 ? dirty_1_140 : _GEN_5799; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6322 = _T_7 ? dirty_1_141 : _GEN_5800; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6323 = _T_7 ? dirty_1_142 : _GEN_5801; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6324 = _T_7 ? dirty_1_143 : _GEN_5802; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6325 = _T_7 ? dirty_1_144 : _GEN_5803; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6326 = _T_7 ? dirty_1_145 : _GEN_5804; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6327 = _T_7 ? dirty_1_146 : _GEN_5805; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6328 = _T_7 ? dirty_1_147 : _GEN_5806; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6329 = _T_7 ? dirty_1_148 : _GEN_5807; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6330 = _T_7 ? dirty_1_149 : _GEN_5808; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6331 = _T_7 ? dirty_1_150 : _GEN_5809; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6332 = _T_7 ? dirty_1_151 : _GEN_5810; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6333 = _T_7 ? dirty_1_152 : _GEN_5811; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6334 = _T_7 ? dirty_1_153 : _GEN_5812; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6335 = _T_7 ? dirty_1_154 : _GEN_5813; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6336 = _T_7 ? dirty_1_155 : _GEN_5814; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6337 = _T_7 ? dirty_1_156 : _GEN_5815; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6338 = _T_7 ? dirty_1_157 : _GEN_5816; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6339 = _T_7 ? dirty_1_158 : _GEN_5817; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6340 = _T_7 ? dirty_1_159 : _GEN_5818; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6341 = _T_7 ? dirty_1_160 : _GEN_5819; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6342 = _T_7 ? dirty_1_161 : _GEN_5820; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6343 = _T_7 ? dirty_1_162 : _GEN_5821; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6344 = _T_7 ? dirty_1_163 : _GEN_5822; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6345 = _T_7 ? dirty_1_164 : _GEN_5823; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6346 = _T_7 ? dirty_1_165 : _GEN_5824; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6347 = _T_7 ? dirty_1_166 : _GEN_5825; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6348 = _T_7 ? dirty_1_167 : _GEN_5826; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6349 = _T_7 ? dirty_1_168 : _GEN_5827; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6350 = _T_7 ? dirty_1_169 : _GEN_5828; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6351 = _T_7 ? dirty_1_170 : _GEN_5829; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6352 = _T_7 ? dirty_1_171 : _GEN_5830; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6353 = _T_7 ? dirty_1_172 : _GEN_5831; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6354 = _T_7 ? dirty_1_173 : _GEN_5832; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6355 = _T_7 ? dirty_1_174 : _GEN_5833; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6356 = _T_7 ? dirty_1_175 : _GEN_5834; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6357 = _T_7 ? dirty_1_176 : _GEN_5835; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6358 = _T_7 ? dirty_1_177 : _GEN_5836; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6359 = _T_7 ? dirty_1_178 : _GEN_5837; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6360 = _T_7 ? dirty_1_179 : _GEN_5838; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6361 = _T_7 ? dirty_1_180 : _GEN_5839; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6362 = _T_7 ? dirty_1_181 : _GEN_5840; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6363 = _T_7 ? dirty_1_182 : _GEN_5841; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6364 = _T_7 ? dirty_1_183 : _GEN_5842; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6365 = _T_7 ? dirty_1_184 : _GEN_5843; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6366 = _T_7 ? dirty_1_185 : _GEN_5844; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6367 = _T_7 ? dirty_1_186 : _GEN_5845; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6368 = _T_7 ? dirty_1_187 : _GEN_5846; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6369 = _T_7 ? dirty_1_188 : _GEN_5847; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6370 = _T_7 ? dirty_1_189 : _GEN_5848; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6371 = _T_7 ? dirty_1_190 : _GEN_5849; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6372 = _T_7 ? dirty_1_191 : _GEN_5850; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6373 = _T_7 ? dirty_1_192 : _GEN_5851; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6374 = _T_7 ? dirty_1_193 : _GEN_5852; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6375 = _T_7 ? dirty_1_194 : _GEN_5853; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6376 = _T_7 ? dirty_1_195 : _GEN_5854; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6377 = _T_7 ? dirty_1_196 : _GEN_5855; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6378 = _T_7 ? dirty_1_197 : _GEN_5856; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6379 = _T_7 ? dirty_1_198 : _GEN_5857; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6380 = _T_7 ? dirty_1_199 : _GEN_5858; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6381 = _T_7 ? dirty_1_200 : _GEN_5859; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6382 = _T_7 ? dirty_1_201 : _GEN_5860; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6383 = _T_7 ? dirty_1_202 : _GEN_5861; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6384 = _T_7 ? dirty_1_203 : _GEN_5862; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6385 = _T_7 ? dirty_1_204 : _GEN_5863; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6386 = _T_7 ? dirty_1_205 : _GEN_5864; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6387 = _T_7 ? dirty_1_206 : _GEN_5865; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6388 = _T_7 ? dirty_1_207 : _GEN_5866; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6389 = _T_7 ? dirty_1_208 : _GEN_5867; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6390 = _T_7 ? dirty_1_209 : _GEN_5868; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6391 = _T_7 ? dirty_1_210 : _GEN_5869; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6392 = _T_7 ? dirty_1_211 : _GEN_5870; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6393 = _T_7 ? dirty_1_212 : _GEN_5871; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6394 = _T_7 ? dirty_1_213 : _GEN_5872; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6395 = _T_7 ? dirty_1_214 : _GEN_5873; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6396 = _T_7 ? dirty_1_215 : _GEN_5874; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6397 = _T_7 ? dirty_1_216 : _GEN_5875; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6398 = _T_7 ? dirty_1_217 : _GEN_5876; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6399 = _T_7 ? dirty_1_218 : _GEN_5877; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6400 = _T_7 ? dirty_1_219 : _GEN_5878; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6401 = _T_7 ? dirty_1_220 : _GEN_5879; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6402 = _T_7 ? dirty_1_221 : _GEN_5880; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6403 = _T_7 ? dirty_1_222 : _GEN_5881; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6404 = _T_7 ? dirty_1_223 : _GEN_5882; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6405 = _T_7 ? dirty_1_224 : _GEN_5883; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6406 = _T_7 ? dirty_1_225 : _GEN_5884; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6407 = _T_7 ? dirty_1_226 : _GEN_5885; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6408 = _T_7 ? dirty_1_227 : _GEN_5886; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6409 = _T_7 ? dirty_1_228 : _GEN_5887; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6410 = _T_7 ? dirty_1_229 : _GEN_5888; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6411 = _T_7 ? dirty_1_230 : _GEN_5889; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6412 = _T_7 ? dirty_1_231 : _GEN_5890; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6413 = _T_7 ? dirty_1_232 : _GEN_5891; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6414 = _T_7 ? dirty_1_233 : _GEN_5892; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6415 = _T_7 ? dirty_1_234 : _GEN_5893; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6416 = _T_7 ? dirty_1_235 : _GEN_5894; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6417 = _T_7 ? dirty_1_236 : _GEN_5895; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6418 = _T_7 ? dirty_1_237 : _GEN_5896; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6419 = _T_7 ? dirty_1_238 : _GEN_5897; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6420 = _T_7 ? dirty_1_239 : _GEN_5898; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6421 = _T_7 ? dirty_1_240 : _GEN_5899; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6422 = _T_7 ? dirty_1_241 : _GEN_5900; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6423 = _T_7 ? dirty_1_242 : _GEN_5901; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6424 = _T_7 ? dirty_1_243 : _GEN_5902; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6425 = _T_7 ? dirty_1_244 : _GEN_5903; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6426 = _T_7 ? dirty_1_245 : _GEN_5904; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6427 = _T_7 ? dirty_1_246 : _GEN_5905; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6428 = _T_7 ? dirty_1_247 : _GEN_5906; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6429 = _T_7 ? dirty_1_248 : _GEN_5907; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6430 = _T_7 ? dirty_1_249 : _GEN_5908; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6431 = _T_7 ? dirty_1_250 : _GEN_5909; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6432 = _T_7 ? dirty_1_251 : _GEN_5910; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6433 = _T_7 ? dirty_1_252 : _GEN_5911; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6434 = _T_7 ? dirty_1_253 : _GEN_5912; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6435 = _T_7 ? dirty_1_254 : _GEN_5913; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6436 = _T_7 ? dirty_1_255 : _GEN_5914; // @[dcache.scala 113:28 397:36]
  wire  _GEN_6437 = _T_7 & cacheInst_r; // @[dcache.scala 397:36 89:38 427:61]
  wire  _GEN_6438 = _T_7 & invalidate; // @[dcache.scala 397:36 90:38 428:61]
  wire  _GEN_6439 = _T_7 & indexOnly; // @[dcache.scala 397:36 94:38 429:61]
  wire  _GEN_6440 = _T_7 & writeBack; // @[dcache.scala 397:36 93:38 430:61]
  wire  _GEN_6441 = _T_7 & storeTag; // @[dcache.scala 397:36 92:38 431:61]
  wire  _GEN_6442 = _T_7 & loadTag; // @[dcache.scala 397:36 91:38 432:61]
  wire [1:0] _GEN_6443 = _T_49 ? _GEN_1766 : wr_cnt; // @[dcache.scala 382:13 178:34]
  wire [31:0] _GEN_6444 = _T_49 ? _GEN_1767 : 32'h0; // @[dcache.scala 382:13 149:33]
  wire [31:0] _GEN_6445 = _T_49 ? _GEN_1768 : 32'h0; // @[dcache.scala 382:13 149:33]
  wire [31:0] _GEN_6446 = _T_49 ? _GEN_1769 : 32'h0; // @[dcache.scala 382:13 149:33]
  wire [31:0] _GEN_6447 = _T_49 ? _GEN_1770 : 32'h0; // @[dcache.scala 382:13 149:33]
  wire [31:0] _GEN_6448 = _T_49 ? _GEN_1771 : 32'h0; // @[dcache.scala 382:13 149:33]
  wire [31:0] _GEN_6449 = _T_49 ? _GEN_1772 : 32'h0; // @[dcache.scala 382:13 149:33]
  wire [31:0] _GEN_6450 = _T_49 ? _GEN_1773 : 32'h0; // @[dcache.scala 382:13 149:33]
  wire [31:0] _GEN_6451 = _T_49 ? _GEN_1774 : 32'h0; // @[dcache.scala 382:13 149:33]
  wire [3:0] _GEN_6452 = _T_49 ? _GEN_1775 : 4'h0; // @[dcache.scala 382:13 150:33]
  wire [3:0] _GEN_6453 = _T_49 ? _GEN_1776 : 4'h0; // @[dcache.scala 382:13 150:33]
  wire [3:0] _GEN_6454 = _T_49 ? _GEN_1777 : 4'h0; // @[dcache.scala 382:13 150:33]
  wire [3:0] _GEN_6455 = _T_49 ? _GEN_1778 : 4'h0; // @[dcache.scala 382:13 150:33]
  wire [3:0] _GEN_6456 = _T_49 ? _GEN_1779 : 4'h0; // @[dcache.scala 382:13 150:33]
  wire [3:0] _GEN_6457 = _T_49 ? _GEN_1780 : 4'h0; // @[dcache.scala 382:13 150:33]
  wire [3:0] _GEN_6458 = _T_49 ? _GEN_1781 : 4'h0; // @[dcache.scala 382:13 150:33]
  wire [3:0] _GEN_6459 = _T_49 ? _GEN_1782 : 4'h0; // @[dcache.scala 382:13 150:33]
  wire [2:0] _GEN_6460 = _T_49 ? _GEN_1783 : _GEN_5917; // @[dcache.scala 382:13]
  wire  _GEN_6461 = _T_49 ? _GEN_1784 : _GEN_5925; // @[dcache.scala 382:13]
  wire  _GEN_6462 = _T_49 ? _GEN_1785 : _GEN_5926; // @[dcache.scala 382:13]
  wire  _GEN_6463 = _T_49 ? _GEN_1786 : _GEN_5927; // @[dcache.scala 382:13]
  wire  _GEN_6464 = _T_49 ? _GEN_1787 : _GEN_5928; // @[dcache.scala 382:13]
  wire  _GEN_6465 = _T_49 ? _GEN_1788 : _GEN_5929; // @[dcache.scala 382:13]
  wire  _GEN_6466 = _T_49 ? _GEN_1789 : _GEN_5930; // @[dcache.scala 382:13]
  wire  _GEN_6467 = _T_49 ? _GEN_1790 : _GEN_5931; // @[dcache.scala 382:13]
  wire  _GEN_6468 = _T_49 ? _GEN_1791 : _GEN_5932; // @[dcache.scala 382:13]
  wire  _GEN_6469 = _T_49 ? _GEN_1792 : _GEN_5933; // @[dcache.scala 382:13]
  wire  _GEN_6470 = _T_49 ? _GEN_1793 : _GEN_5934; // @[dcache.scala 382:13]
  wire  _GEN_6471 = _T_49 ? _GEN_1794 : _GEN_5935; // @[dcache.scala 382:13]
  wire  _GEN_6472 = _T_49 ? _GEN_1795 : _GEN_5936; // @[dcache.scala 382:13]
  wire  _GEN_6473 = _T_49 ? _GEN_1796 : _GEN_5937; // @[dcache.scala 382:13]
  wire  _GEN_6474 = _T_49 ? _GEN_1797 : _GEN_5938; // @[dcache.scala 382:13]
  wire  _GEN_6475 = _T_49 ? _GEN_1798 : _GEN_5939; // @[dcache.scala 382:13]
  wire  _GEN_6476 = _T_49 ? _GEN_1799 : _GEN_5940; // @[dcache.scala 382:13]
  wire  _GEN_6477 = _T_49 ? _GEN_1800 : _GEN_5941; // @[dcache.scala 382:13]
  wire  _GEN_6478 = _T_49 ? _GEN_1801 : _GEN_5942; // @[dcache.scala 382:13]
  wire  _GEN_6479 = _T_49 ? _GEN_1802 : _GEN_5943; // @[dcache.scala 382:13]
  wire  _GEN_6480 = _T_49 ? _GEN_1803 : _GEN_5944; // @[dcache.scala 382:13]
  wire  _GEN_6481 = _T_49 ? _GEN_1804 : _GEN_5945; // @[dcache.scala 382:13]
  wire  _GEN_6482 = _T_49 ? _GEN_1805 : _GEN_5946; // @[dcache.scala 382:13]
  wire  _GEN_6483 = _T_49 ? _GEN_1806 : _GEN_5947; // @[dcache.scala 382:13]
  wire  _GEN_6484 = _T_49 ? _GEN_1807 : _GEN_5948; // @[dcache.scala 382:13]
  wire  _GEN_6485 = _T_49 ? _GEN_1808 : _GEN_5949; // @[dcache.scala 382:13]
  wire  _GEN_6486 = _T_49 ? _GEN_1809 : _GEN_5950; // @[dcache.scala 382:13]
  wire  _GEN_6487 = _T_49 ? _GEN_1810 : _GEN_5951; // @[dcache.scala 382:13]
  wire  _GEN_6488 = _T_49 ? _GEN_1811 : _GEN_5952; // @[dcache.scala 382:13]
  wire  _GEN_6489 = _T_49 ? _GEN_1812 : _GEN_5953; // @[dcache.scala 382:13]
  wire  _GEN_6490 = _T_49 ? _GEN_1813 : _GEN_5954; // @[dcache.scala 382:13]
  wire  _GEN_6491 = _T_49 ? _GEN_1814 : _GEN_5955; // @[dcache.scala 382:13]
  wire  _GEN_6492 = _T_49 ? _GEN_1815 : _GEN_5956; // @[dcache.scala 382:13]
  wire  _GEN_6493 = _T_49 ? _GEN_1816 : _GEN_5957; // @[dcache.scala 382:13]
  wire  _GEN_6494 = _T_49 ? _GEN_1817 : _GEN_5958; // @[dcache.scala 382:13]
  wire  _GEN_6495 = _T_49 ? _GEN_1818 : _GEN_5959; // @[dcache.scala 382:13]
  wire  _GEN_6496 = _T_49 ? _GEN_1819 : _GEN_5960; // @[dcache.scala 382:13]
  wire  _GEN_6497 = _T_49 ? _GEN_1820 : _GEN_5961; // @[dcache.scala 382:13]
  wire  _GEN_6498 = _T_49 ? _GEN_1821 : _GEN_5962; // @[dcache.scala 382:13]
  wire  _GEN_6499 = _T_49 ? _GEN_1822 : _GEN_5963; // @[dcache.scala 382:13]
  wire  _GEN_6500 = _T_49 ? _GEN_1823 : _GEN_5964; // @[dcache.scala 382:13]
  wire  _GEN_6501 = _T_49 ? _GEN_1824 : _GEN_5965; // @[dcache.scala 382:13]
  wire  _GEN_6502 = _T_49 ? _GEN_1825 : _GEN_5966; // @[dcache.scala 382:13]
  wire  _GEN_6503 = _T_49 ? _GEN_1826 : _GEN_5967; // @[dcache.scala 382:13]
  wire  _GEN_6504 = _T_49 ? _GEN_1827 : _GEN_5968; // @[dcache.scala 382:13]
  wire  _GEN_6505 = _T_49 ? _GEN_1828 : _GEN_5969; // @[dcache.scala 382:13]
  wire  _GEN_6506 = _T_49 ? _GEN_1829 : _GEN_5970; // @[dcache.scala 382:13]
  wire  _GEN_6507 = _T_49 ? _GEN_1830 : _GEN_5971; // @[dcache.scala 382:13]
  wire  _GEN_6508 = _T_49 ? _GEN_1831 : _GEN_5972; // @[dcache.scala 382:13]
  wire  _GEN_6509 = _T_49 ? _GEN_1832 : _GEN_5973; // @[dcache.scala 382:13]
  wire  _GEN_6510 = _T_49 ? _GEN_1833 : _GEN_5974; // @[dcache.scala 382:13]
  wire  _GEN_6511 = _T_49 ? _GEN_1834 : _GEN_5975; // @[dcache.scala 382:13]
  wire  _GEN_6512 = _T_49 ? _GEN_1835 : _GEN_5976; // @[dcache.scala 382:13]
  wire  _GEN_6513 = _T_49 ? _GEN_1836 : _GEN_5977; // @[dcache.scala 382:13]
  wire  _GEN_6514 = _T_49 ? _GEN_1837 : _GEN_5978; // @[dcache.scala 382:13]
  wire  _GEN_6515 = _T_49 ? _GEN_1838 : _GEN_5979; // @[dcache.scala 382:13]
  wire  _GEN_6516 = _T_49 ? _GEN_1839 : _GEN_5980; // @[dcache.scala 382:13]
  wire  _GEN_6517 = _T_49 ? _GEN_1840 : _GEN_5981; // @[dcache.scala 382:13]
  wire  _GEN_6518 = _T_49 ? _GEN_1841 : _GEN_5982; // @[dcache.scala 382:13]
  wire  _GEN_6519 = _T_49 ? _GEN_1842 : _GEN_5983; // @[dcache.scala 382:13]
  wire  _GEN_6520 = _T_49 ? _GEN_1843 : _GEN_5984; // @[dcache.scala 382:13]
  wire  _GEN_6521 = _T_49 ? _GEN_1844 : _GEN_5985; // @[dcache.scala 382:13]
  wire  _GEN_6522 = _T_49 ? _GEN_1845 : _GEN_5986; // @[dcache.scala 382:13]
  wire  _GEN_6523 = _T_49 ? _GEN_1846 : _GEN_5987; // @[dcache.scala 382:13]
  wire  _GEN_6524 = _T_49 ? _GEN_1847 : _GEN_5988; // @[dcache.scala 382:13]
  wire  _GEN_6525 = _T_49 ? _GEN_1848 : _GEN_5989; // @[dcache.scala 382:13]
  wire  _GEN_6526 = _T_49 ? _GEN_1849 : _GEN_5990; // @[dcache.scala 382:13]
  wire  _GEN_6527 = _T_49 ? _GEN_1850 : _GEN_5991; // @[dcache.scala 382:13]
  wire  _GEN_6528 = _T_49 ? _GEN_1851 : _GEN_5992; // @[dcache.scala 382:13]
  wire  _GEN_6529 = _T_49 ? _GEN_1852 : _GEN_5993; // @[dcache.scala 382:13]
  wire  _GEN_6530 = _T_49 ? _GEN_1853 : _GEN_5994; // @[dcache.scala 382:13]
  wire  _GEN_6531 = _T_49 ? _GEN_1854 : _GEN_5995; // @[dcache.scala 382:13]
  wire  _GEN_6532 = _T_49 ? _GEN_1855 : _GEN_5996; // @[dcache.scala 382:13]
  wire  _GEN_6533 = _T_49 ? _GEN_1856 : _GEN_5997; // @[dcache.scala 382:13]
  wire  _GEN_6534 = _T_49 ? _GEN_1857 : _GEN_5998; // @[dcache.scala 382:13]
  wire  _GEN_6535 = _T_49 ? _GEN_1858 : _GEN_5999; // @[dcache.scala 382:13]
  wire  _GEN_6536 = _T_49 ? _GEN_1859 : _GEN_6000; // @[dcache.scala 382:13]
  wire  _GEN_6537 = _T_49 ? _GEN_1860 : _GEN_6001; // @[dcache.scala 382:13]
  wire  _GEN_6538 = _T_49 ? _GEN_1861 : _GEN_6002; // @[dcache.scala 382:13]
  wire  _GEN_6539 = _T_49 ? _GEN_1862 : _GEN_6003; // @[dcache.scala 382:13]
  wire  _GEN_6540 = _T_49 ? _GEN_1863 : _GEN_6004; // @[dcache.scala 382:13]
  wire  _GEN_6541 = _T_49 ? _GEN_1864 : _GEN_6005; // @[dcache.scala 382:13]
  wire  _GEN_6542 = _T_49 ? _GEN_1865 : _GEN_6006; // @[dcache.scala 382:13]
  wire  _GEN_6543 = _T_49 ? _GEN_1866 : _GEN_6007; // @[dcache.scala 382:13]
  wire  _GEN_6544 = _T_49 ? _GEN_1867 : _GEN_6008; // @[dcache.scala 382:13]
  wire  _GEN_6545 = _T_49 ? _GEN_1868 : _GEN_6009; // @[dcache.scala 382:13]
  wire  _GEN_6546 = _T_49 ? _GEN_1869 : _GEN_6010; // @[dcache.scala 382:13]
  wire  _GEN_6547 = _T_49 ? _GEN_1870 : _GEN_6011; // @[dcache.scala 382:13]
  wire  _GEN_6548 = _T_49 ? _GEN_1871 : _GEN_6012; // @[dcache.scala 382:13]
  wire  _GEN_6549 = _T_49 ? _GEN_1872 : _GEN_6013; // @[dcache.scala 382:13]
  wire  _GEN_6550 = _T_49 ? _GEN_1873 : _GEN_6014; // @[dcache.scala 382:13]
  wire  _GEN_6551 = _T_49 ? _GEN_1874 : _GEN_6015; // @[dcache.scala 382:13]
  wire  _GEN_6552 = _T_49 ? _GEN_1875 : _GEN_6016; // @[dcache.scala 382:13]
  wire  _GEN_6553 = _T_49 ? _GEN_1876 : _GEN_6017; // @[dcache.scala 382:13]
  wire  _GEN_6554 = _T_49 ? _GEN_1877 : _GEN_6018; // @[dcache.scala 382:13]
  wire  _GEN_6555 = _T_49 ? _GEN_1878 : _GEN_6019; // @[dcache.scala 382:13]
  wire  _GEN_6556 = _T_49 ? _GEN_1879 : _GEN_6020; // @[dcache.scala 382:13]
  wire  _GEN_6557 = _T_49 ? _GEN_1880 : _GEN_6021; // @[dcache.scala 382:13]
  wire  _GEN_6558 = _T_49 ? _GEN_1881 : _GEN_6022; // @[dcache.scala 382:13]
  wire  _GEN_6559 = _T_49 ? _GEN_1882 : _GEN_6023; // @[dcache.scala 382:13]
  wire  _GEN_6560 = _T_49 ? _GEN_1883 : _GEN_6024; // @[dcache.scala 382:13]
  wire  _GEN_6561 = _T_49 ? _GEN_1884 : _GEN_6025; // @[dcache.scala 382:13]
  wire  _GEN_6562 = _T_49 ? _GEN_1885 : _GEN_6026; // @[dcache.scala 382:13]
  wire  _GEN_6563 = _T_49 ? _GEN_1886 : _GEN_6027; // @[dcache.scala 382:13]
  wire  _GEN_6564 = _T_49 ? _GEN_1887 : _GEN_6028; // @[dcache.scala 382:13]
  wire  _GEN_6565 = _T_49 ? _GEN_1888 : _GEN_6029; // @[dcache.scala 382:13]
  wire  _GEN_6566 = _T_49 ? _GEN_1889 : _GEN_6030; // @[dcache.scala 382:13]
  wire  _GEN_6567 = _T_49 ? _GEN_1890 : _GEN_6031; // @[dcache.scala 382:13]
  wire  _GEN_6568 = _T_49 ? _GEN_1891 : _GEN_6032; // @[dcache.scala 382:13]
  wire  _GEN_6569 = _T_49 ? _GEN_1892 : _GEN_6033; // @[dcache.scala 382:13]
  wire  _GEN_6570 = _T_49 ? _GEN_1893 : _GEN_6034; // @[dcache.scala 382:13]
  wire  _GEN_6571 = _T_49 ? _GEN_1894 : _GEN_6035; // @[dcache.scala 382:13]
  wire  _GEN_6572 = _T_49 ? _GEN_1895 : _GEN_6036; // @[dcache.scala 382:13]
  wire  _GEN_6573 = _T_49 ? _GEN_1896 : _GEN_6037; // @[dcache.scala 382:13]
  wire  _GEN_6574 = _T_49 ? _GEN_1897 : _GEN_6038; // @[dcache.scala 382:13]
  wire  _GEN_6575 = _T_49 ? _GEN_1898 : _GEN_6039; // @[dcache.scala 382:13]
  wire  _GEN_6576 = _T_49 ? _GEN_1899 : _GEN_6040; // @[dcache.scala 382:13]
  wire  _GEN_6577 = _T_49 ? _GEN_1900 : _GEN_6041; // @[dcache.scala 382:13]
  wire  _GEN_6578 = _T_49 ? _GEN_1901 : _GEN_6042; // @[dcache.scala 382:13]
  wire  _GEN_6579 = _T_49 ? _GEN_1902 : _GEN_6043; // @[dcache.scala 382:13]
  wire  _GEN_6580 = _T_49 ? _GEN_1903 : _GEN_6044; // @[dcache.scala 382:13]
  wire  _GEN_6581 = _T_49 ? _GEN_1904 : _GEN_6045; // @[dcache.scala 382:13]
  wire  _GEN_6582 = _T_49 ? _GEN_1905 : _GEN_6046; // @[dcache.scala 382:13]
  wire  _GEN_6583 = _T_49 ? _GEN_1906 : _GEN_6047; // @[dcache.scala 382:13]
  wire  _GEN_6584 = _T_49 ? _GEN_1907 : _GEN_6048; // @[dcache.scala 382:13]
  wire  _GEN_6585 = _T_49 ? _GEN_1908 : _GEN_6049; // @[dcache.scala 382:13]
  wire  _GEN_6586 = _T_49 ? _GEN_1909 : _GEN_6050; // @[dcache.scala 382:13]
  wire  _GEN_6587 = _T_49 ? _GEN_1910 : _GEN_6051; // @[dcache.scala 382:13]
  wire  _GEN_6588 = _T_49 ? _GEN_1911 : _GEN_6052; // @[dcache.scala 382:13]
  wire  _GEN_6589 = _T_49 ? _GEN_1912 : _GEN_6053; // @[dcache.scala 382:13]
  wire  _GEN_6590 = _T_49 ? _GEN_1913 : _GEN_6054; // @[dcache.scala 382:13]
  wire  _GEN_6591 = _T_49 ? _GEN_1914 : _GEN_6055; // @[dcache.scala 382:13]
  wire  _GEN_6592 = _T_49 ? _GEN_1915 : _GEN_6056; // @[dcache.scala 382:13]
  wire  _GEN_6593 = _T_49 ? _GEN_1916 : _GEN_6057; // @[dcache.scala 382:13]
  wire  _GEN_6594 = _T_49 ? _GEN_1917 : _GEN_6058; // @[dcache.scala 382:13]
  wire  _GEN_6595 = _T_49 ? _GEN_1918 : _GEN_6059; // @[dcache.scala 382:13]
  wire  _GEN_6596 = _T_49 ? _GEN_1919 : _GEN_6060; // @[dcache.scala 382:13]
  wire  _GEN_6597 = _T_49 ? _GEN_1920 : _GEN_6061; // @[dcache.scala 382:13]
  wire  _GEN_6598 = _T_49 ? _GEN_1921 : _GEN_6062; // @[dcache.scala 382:13]
  wire  _GEN_6599 = _T_49 ? _GEN_1922 : _GEN_6063; // @[dcache.scala 382:13]
  wire  _GEN_6600 = _T_49 ? _GEN_1923 : _GEN_6064; // @[dcache.scala 382:13]
  wire  _GEN_6601 = _T_49 ? _GEN_1924 : _GEN_6065; // @[dcache.scala 382:13]
  wire  _GEN_6602 = _T_49 ? _GEN_1925 : _GEN_6066; // @[dcache.scala 382:13]
  wire  _GEN_6603 = _T_49 ? _GEN_1926 : _GEN_6067; // @[dcache.scala 382:13]
  wire  _GEN_6604 = _T_49 ? _GEN_1927 : _GEN_6068; // @[dcache.scala 382:13]
  wire  _GEN_6605 = _T_49 ? _GEN_1928 : _GEN_6069; // @[dcache.scala 382:13]
  wire  _GEN_6606 = _T_49 ? _GEN_1929 : _GEN_6070; // @[dcache.scala 382:13]
  wire  _GEN_6607 = _T_49 ? _GEN_1930 : _GEN_6071; // @[dcache.scala 382:13]
  wire  _GEN_6608 = _T_49 ? _GEN_1931 : _GEN_6072; // @[dcache.scala 382:13]
  wire  _GEN_6609 = _T_49 ? _GEN_1932 : _GEN_6073; // @[dcache.scala 382:13]
  wire  _GEN_6610 = _T_49 ? _GEN_1933 : _GEN_6074; // @[dcache.scala 382:13]
  wire  _GEN_6611 = _T_49 ? _GEN_1934 : _GEN_6075; // @[dcache.scala 382:13]
  wire  _GEN_6612 = _T_49 ? _GEN_1935 : _GEN_6076; // @[dcache.scala 382:13]
  wire  _GEN_6613 = _T_49 ? _GEN_1936 : _GEN_6077; // @[dcache.scala 382:13]
  wire  _GEN_6614 = _T_49 ? _GEN_1937 : _GEN_6078; // @[dcache.scala 382:13]
  wire  _GEN_6615 = _T_49 ? _GEN_1938 : _GEN_6079; // @[dcache.scala 382:13]
  wire  _GEN_6616 = _T_49 ? _GEN_1939 : _GEN_6080; // @[dcache.scala 382:13]
  wire  _GEN_6617 = _T_49 ? _GEN_1940 : _GEN_6081; // @[dcache.scala 382:13]
  wire  _GEN_6618 = _T_49 ? _GEN_1941 : _GEN_6082; // @[dcache.scala 382:13]
  wire  _GEN_6619 = _T_49 ? _GEN_1942 : _GEN_6083; // @[dcache.scala 382:13]
  wire  _GEN_6620 = _T_49 ? _GEN_1943 : _GEN_6084; // @[dcache.scala 382:13]
  wire  _GEN_6621 = _T_49 ? _GEN_1944 : _GEN_6085; // @[dcache.scala 382:13]
  wire  _GEN_6622 = _T_49 ? _GEN_1945 : _GEN_6086; // @[dcache.scala 382:13]
  wire  _GEN_6623 = _T_49 ? _GEN_1946 : _GEN_6087; // @[dcache.scala 382:13]
  wire  _GEN_6624 = _T_49 ? _GEN_1947 : _GEN_6088; // @[dcache.scala 382:13]
  wire  _GEN_6625 = _T_49 ? _GEN_1948 : _GEN_6089; // @[dcache.scala 382:13]
  wire  _GEN_6626 = _T_49 ? _GEN_1949 : _GEN_6090; // @[dcache.scala 382:13]
  wire  _GEN_6627 = _T_49 ? _GEN_1950 : _GEN_6091; // @[dcache.scala 382:13]
  wire  _GEN_6628 = _T_49 ? _GEN_1951 : _GEN_6092; // @[dcache.scala 382:13]
  wire  _GEN_6629 = _T_49 ? _GEN_1952 : _GEN_6093; // @[dcache.scala 382:13]
  wire  _GEN_6630 = _T_49 ? _GEN_1953 : _GEN_6094; // @[dcache.scala 382:13]
  wire  _GEN_6631 = _T_49 ? _GEN_1954 : _GEN_6095; // @[dcache.scala 382:13]
  wire  _GEN_6632 = _T_49 ? _GEN_1955 : _GEN_6096; // @[dcache.scala 382:13]
  wire  _GEN_6633 = _T_49 ? _GEN_1956 : _GEN_6097; // @[dcache.scala 382:13]
  wire  _GEN_6634 = _T_49 ? _GEN_1957 : _GEN_6098; // @[dcache.scala 382:13]
  wire  _GEN_6635 = _T_49 ? _GEN_1958 : _GEN_6099; // @[dcache.scala 382:13]
  wire  _GEN_6636 = _T_49 ? _GEN_1959 : _GEN_6100; // @[dcache.scala 382:13]
  wire  _GEN_6637 = _T_49 ? _GEN_1960 : _GEN_6101; // @[dcache.scala 382:13]
  wire  _GEN_6638 = _T_49 ? _GEN_1961 : _GEN_6102; // @[dcache.scala 382:13]
  wire  _GEN_6639 = _T_49 ? _GEN_1962 : _GEN_6103; // @[dcache.scala 382:13]
  wire  _GEN_6640 = _T_49 ? _GEN_1963 : _GEN_6104; // @[dcache.scala 382:13]
  wire  _GEN_6641 = _T_49 ? _GEN_1964 : _GEN_6105; // @[dcache.scala 382:13]
  wire  _GEN_6642 = _T_49 ? _GEN_1965 : _GEN_6106; // @[dcache.scala 382:13]
  wire  _GEN_6643 = _T_49 ? _GEN_1966 : _GEN_6107; // @[dcache.scala 382:13]
  wire  _GEN_6644 = _T_49 ? _GEN_1967 : _GEN_6108; // @[dcache.scala 382:13]
  wire  _GEN_6645 = _T_49 ? _GEN_1968 : _GEN_6109; // @[dcache.scala 382:13]
  wire  _GEN_6646 = _T_49 ? _GEN_1969 : _GEN_6110; // @[dcache.scala 382:13]
  wire  _GEN_6647 = _T_49 ? _GEN_1970 : _GEN_6111; // @[dcache.scala 382:13]
  wire  _GEN_6648 = _T_49 ? _GEN_1971 : _GEN_6112; // @[dcache.scala 382:13]
  wire  _GEN_6649 = _T_49 ? _GEN_1972 : _GEN_6113; // @[dcache.scala 382:13]
  wire  _GEN_6650 = _T_49 ? _GEN_1973 : _GEN_6114; // @[dcache.scala 382:13]
  wire  _GEN_6651 = _T_49 ? _GEN_1974 : _GEN_6115; // @[dcache.scala 382:13]
  wire  _GEN_6652 = _T_49 ? _GEN_1975 : _GEN_6116; // @[dcache.scala 382:13]
  wire  _GEN_6653 = _T_49 ? _GEN_1976 : _GEN_6117; // @[dcache.scala 382:13]
  wire  _GEN_6654 = _T_49 ? _GEN_1977 : _GEN_6118; // @[dcache.scala 382:13]
  wire  _GEN_6655 = _T_49 ? _GEN_1978 : _GEN_6119; // @[dcache.scala 382:13]
  wire  _GEN_6656 = _T_49 ? _GEN_1979 : _GEN_6120; // @[dcache.scala 382:13]
  wire  _GEN_6657 = _T_49 ? _GEN_1980 : _GEN_6121; // @[dcache.scala 382:13]
  wire  _GEN_6658 = _T_49 ? _GEN_1981 : _GEN_6122; // @[dcache.scala 382:13]
  wire  _GEN_6659 = _T_49 ? _GEN_1982 : _GEN_6123; // @[dcache.scala 382:13]
  wire  _GEN_6660 = _T_49 ? _GEN_1983 : _GEN_6124; // @[dcache.scala 382:13]
  wire  _GEN_6661 = _T_49 ? _GEN_1984 : _GEN_6125; // @[dcache.scala 382:13]
  wire  _GEN_6662 = _T_49 ? _GEN_1985 : _GEN_6126; // @[dcache.scala 382:13]
  wire  _GEN_6663 = _T_49 ? _GEN_1986 : _GEN_6127; // @[dcache.scala 382:13]
  wire  _GEN_6664 = _T_49 ? _GEN_1987 : _GEN_6128; // @[dcache.scala 382:13]
  wire  _GEN_6665 = _T_49 ? _GEN_1988 : _GEN_6129; // @[dcache.scala 382:13]
  wire  _GEN_6666 = _T_49 ? _GEN_1989 : _GEN_6130; // @[dcache.scala 382:13]
  wire  _GEN_6667 = _T_49 ? _GEN_1990 : _GEN_6131; // @[dcache.scala 382:13]
  wire  _GEN_6668 = _T_49 ? _GEN_1991 : _GEN_6132; // @[dcache.scala 382:13]
  wire  _GEN_6669 = _T_49 ? _GEN_1992 : _GEN_6133; // @[dcache.scala 382:13]
  wire  _GEN_6670 = _T_49 ? _GEN_1993 : _GEN_6134; // @[dcache.scala 382:13]
  wire  _GEN_6671 = _T_49 ? _GEN_1994 : _GEN_6135; // @[dcache.scala 382:13]
  wire  _GEN_6672 = _T_49 ? _GEN_1995 : _GEN_6136; // @[dcache.scala 382:13]
  wire  _GEN_6673 = _T_49 ? _GEN_1996 : _GEN_6137; // @[dcache.scala 382:13]
  wire  _GEN_6674 = _T_49 ? _GEN_1997 : _GEN_6138; // @[dcache.scala 382:13]
  wire  _GEN_6675 = _T_49 ? _GEN_1998 : _GEN_6139; // @[dcache.scala 382:13]
  wire  _GEN_6676 = _T_49 ? _GEN_1999 : _GEN_6140; // @[dcache.scala 382:13]
  wire  _GEN_6677 = _T_49 ? _GEN_2000 : _GEN_6141; // @[dcache.scala 382:13]
  wire  _GEN_6678 = _T_49 ? _GEN_2001 : _GEN_6142; // @[dcache.scala 382:13]
  wire  _GEN_6679 = _T_49 ? _GEN_2002 : _GEN_6143; // @[dcache.scala 382:13]
  wire  _GEN_6680 = _T_49 ? _GEN_2003 : _GEN_6144; // @[dcache.scala 382:13]
  wire  _GEN_6681 = _T_49 ? _GEN_2004 : _GEN_6145; // @[dcache.scala 382:13]
  wire  _GEN_6682 = _T_49 ? _GEN_2005 : _GEN_6146; // @[dcache.scala 382:13]
  wire  _GEN_6683 = _T_49 ? _GEN_2006 : _GEN_6147; // @[dcache.scala 382:13]
  wire  _GEN_6684 = _T_49 ? _GEN_2007 : _GEN_6148; // @[dcache.scala 382:13]
  wire  _GEN_6685 = _T_49 ? _GEN_2008 : _GEN_6149; // @[dcache.scala 382:13]
  wire  _GEN_6686 = _T_49 ? _GEN_2009 : _GEN_6150; // @[dcache.scala 382:13]
  wire  _GEN_6687 = _T_49 ? _GEN_2010 : _GEN_6151; // @[dcache.scala 382:13]
  wire  _GEN_6688 = _T_49 ? _GEN_2011 : _GEN_6152; // @[dcache.scala 382:13]
  wire  _GEN_6689 = _T_49 ? _GEN_2012 : _GEN_6153; // @[dcache.scala 382:13]
  wire  _GEN_6690 = _T_49 ? _GEN_2013 : _GEN_6154; // @[dcache.scala 382:13]
  wire  _GEN_6691 = _T_49 ? _GEN_2014 : _GEN_6155; // @[dcache.scala 382:13]
  wire  _GEN_6692 = _T_49 ? _GEN_2015 : _GEN_6156; // @[dcache.scala 382:13]
  wire  _GEN_6693 = _T_49 ? _GEN_2016 : _GEN_6157; // @[dcache.scala 382:13]
  wire  _GEN_6694 = _T_49 ? _GEN_2017 : _GEN_6158; // @[dcache.scala 382:13]
  wire  _GEN_6695 = _T_49 ? _GEN_2018 : _GEN_6159; // @[dcache.scala 382:13]
  wire  _GEN_6696 = _T_49 ? _GEN_2019 : _GEN_6160; // @[dcache.scala 382:13]
  wire  _GEN_6697 = _T_49 ? _GEN_2020 : _GEN_6161; // @[dcache.scala 382:13]
  wire  _GEN_6698 = _T_49 ? _GEN_2021 : _GEN_6162; // @[dcache.scala 382:13]
  wire  _GEN_6699 = _T_49 ? _GEN_2022 : _GEN_6163; // @[dcache.scala 382:13]
  wire  _GEN_6700 = _T_49 ? _GEN_2023 : _GEN_6164; // @[dcache.scala 382:13]
  wire  _GEN_6701 = _T_49 ? _GEN_2024 : _GEN_6165; // @[dcache.scala 382:13]
  wire  _GEN_6702 = _T_49 ? _GEN_2025 : _GEN_6166; // @[dcache.scala 382:13]
  wire  _GEN_6703 = _T_49 ? _GEN_2026 : _GEN_6167; // @[dcache.scala 382:13]
  wire  _GEN_6704 = _T_49 ? _GEN_2027 : _GEN_6168; // @[dcache.scala 382:13]
  wire  _GEN_6705 = _T_49 ? _GEN_2028 : _GEN_6169; // @[dcache.scala 382:13]
  wire  _GEN_6706 = _T_49 ? _GEN_2029 : _GEN_6170; // @[dcache.scala 382:13]
  wire  _GEN_6707 = _T_49 ? _GEN_2030 : _GEN_6171; // @[dcache.scala 382:13]
  wire  _GEN_6708 = _T_49 ? _GEN_2031 : _GEN_6172; // @[dcache.scala 382:13]
  wire  _GEN_6709 = _T_49 ? _GEN_2032 : _GEN_6173; // @[dcache.scala 382:13]
  wire  _GEN_6710 = _T_49 ? _GEN_2033 : _GEN_6174; // @[dcache.scala 382:13]
  wire  _GEN_6711 = _T_49 ? _GEN_2034 : _GEN_6175; // @[dcache.scala 382:13]
  wire  _GEN_6712 = _T_49 ? _GEN_2035 : _GEN_6176; // @[dcache.scala 382:13]
  wire  _GEN_6713 = _T_49 ? _GEN_2036 : _GEN_6177; // @[dcache.scala 382:13]
  wire  _GEN_6714 = _T_49 ? _GEN_2037 : _GEN_6178; // @[dcache.scala 382:13]
  wire  _GEN_6715 = _T_49 ? _GEN_2038 : _GEN_6179; // @[dcache.scala 382:13]
  wire  _GEN_6716 = _T_49 ? _GEN_2039 : _GEN_6180; // @[dcache.scala 382:13]
  wire  _GEN_6717 = _T_49 ? _GEN_2040 : _GEN_6181; // @[dcache.scala 382:13]
  wire  _GEN_6718 = _T_49 ? _GEN_2041 : _GEN_6182; // @[dcache.scala 382:13]
  wire  _GEN_6719 = _T_49 ? _GEN_2042 : _GEN_6183; // @[dcache.scala 382:13]
  wire  _GEN_6720 = _T_49 ? _GEN_2043 : _GEN_6184; // @[dcache.scala 382:13]
  wire  _GEN_6721 = _T_49 ? _GEN_2044 : _GEN_6185; // @[dcache.scala 382:13]
  wire  _GEN_6722 = _T_49 ? _GEN_2045 : _GEN_6186; // @[dcache.scala 382:13]
  wire  _GEN_6723 = _T_49 ? _GEN_2046 : _GEN_6187; // @[dcache.scala 382:13]
  wire  _GEN_6724 = _T_49 ? _GEN_2047 : _GEN_6188; // @[dcache.scala 382:13]
  wire  _GEN_6725 = _T_49 ? _GEN_2048 : _GEN_6189; // @[dcache.scala 382:13]
  wire  _GEN_6726 = _T_49 ? _GEN_2049 : _GEN_6190; // @[dcache.scala 382:13]
  wire  _GEN_6727 = _T_49 ? _GEN_2050 : _GEN_6191; // @[dcache.scala 382:13]
  wire  _GEN_6728 = _T_49 ? _GEN_2051 : _GEN_6192; // @[dcache.scala 382:13]
  wire  _GEN_6729 = _T_49 ? _GEN_2052 : _GEN_6193; // @[dcache.scala 382:13]
  wire  _GEN_6730 = _T_49 ? _GEN_2053 : _GEN_6194; // @[dcache.scala 382:13]
  wire  _GEN_6731 = _T_49 ? _GEN_2054 : _GEN_6195; // @[dcache.scala 382:13]
  wire  _GEN_6732 = _T_49 ? _GEN_2055 : _GEN_6196; // @[dcache.scala 382:13]
  wire  _GEN_6733 = _T_49 ? _GEN_2056 : _GEN_6197; // @[dcache.scala 382:13]
  wire  _GEN_6734 = _T_49 ? _GEN_2057 : _GEN_6198; // @[dcache.scala 382:13]
  wire  _GEN_6735 = _T_49 ? _GEN_2058 : _GEN_6199; // @[dcache.scala 382:13]
  wire  _GEN_6736 = _T_49 ? _GEN_2059 : _GEN_6200; // @[dcache.scala 382:13]
  wire  _GEN_6737 = _T_49 ? _GEN_2060 : _GEN_6201; // @[dcache.scala 382:13]
  wire  _GEN_6738 = _T_49 ? _GEN_2061 : _GEN_6202; // @[dcache.scala 382:13]
  wire  _GEN_6739 = _T_49 ? _GEN_2062 : _GEN_6203; // @[dcache.scala 382:13]
  wire  _GEN_6740 = _T_49 ? _GEN_2063 : _GEN_6204; // @[dcache.scala 382:13]
  wire  _GEN_6741 = _T_49 ? _GEN_2064 : _GEN_6205; // @[dcache.scala 382:13]
  wire  _GEN_6742 = _T_49 ? _GEN_2065 : _GEN_6206; // @[dcache.scala 382:13]
  wire  _GEN_6743 = _T_49 ? _GEN_2066 : _GEN_6207; // @[dcache.scala 382:13]
  wire  _GEN_6744 = _T_49 ? _GEN_2067 : _GEN_6208; // @[dcache.scala 382:13]
  wire  _GEN_6745 = _T_49 ? _GEN_2068 : _GEN_6209; // @[dcache.scala 382:13]
  wire  _GEN_6746 = _T_49 ? _GEN_2069 : _GEN_6210; // @[dcache.scala 382:13]
  wire  _GEN_6747 = _T_49 ? _GEN_2070 : _GEN_6211; // @[dcache.scala 382:13]
  wire  _GEN_6748 = _T_49 ? _GEN_2071 : _GEN_6212; // @[dcache.scala 382:13]
  wire  _GEN_6749 = _T_49 ? _GEN_2072 : _GEN_6213; // @[dcache.scala 382:13]
  wire  _GEN_6750 = _T_49 ? _GEN_2073 : _GEN_6214; // @[dcache.scala 382:13]
  wire  _GEN_6751 = _T_49 ? _GEN_2074 : _GEN_6215; // @[dcache.scala 382:13]
  wire  _GEN_6752 = _T_49 ? _GEN_2075 : _GEN_6216; // @[dcache.scala 382:13]
  wire  _GEN_6753 = _T_49 ? _GEN_2076 : _GEN_6217; // @[dcache.scala 382:13]
  wire  _GEN_6754 = _T_49 ? _GEN_2077 : _GEN_6218; // @[dcache.scala 382:13]
  wire  _GEN_6755 = _T_49 ? _GEN_2078 : _GEN_6219; // @[dcache.scala 382:13]
  wire  _GEN_6756 = _T_49 ? _GEN_2079 : _GEN_6220; // @[dcache.scala 382:13]
  wire  _GEN_6757 = _T_49 ? _GEN_2080 : _GEN_6221; // @[dcache.scala 382:13]
  wire  _GEN_6758 = _T_49 ? _GEN_2081 : _GEN_6222; // @[dcache.scala 382:13]
  wire  _GEN_6759 = _T_49 ? _GEN_2082 : _GEN_6223; // @[dcache.scala 382:13]
  wire  _GEN_6760 = _T_49 ? _GEN_2083 : _GEN_6224; // @[dcache.scala 382:13]
  wire  _GEN_6761 = _T_49 ? _GEN_2084 : _GEN_6225; // @[dcache.scala 382:13]
  wire  _GEN_6762 = _T_49 ? _GEN_2085 : _GEN_6226; // @[dcache.scala 382:13]
  wire  _GEN_6763 = _T_49 ? _GEN_2086 : _GEN_6227; // @[dcache.scala 382:13]
  wire  _GEN_6764 = _T_49 ? _GEN_2087 : _GEN_6228; // @[dcache.scala 382:13]
  wire  _GEN_6765 = _T_49 ? _GEN_2088 : _GEN_6229; // @[dcache.scala 382:13]
  wire  _GEN_6766 = _T_49 ? _GEN_2089 : _GEN_6230; // @[dcache.scala 382:13]
  wire  _GEN_6767 = _T_49 ? _GEN_2090 : _GEN_6231; // @[dcache.scala 382:13]
  wire  _GEN_6768 = _T_49 ? _GEN_2091 : _GEN_6232; // @[dcache.scala 382:13]
  wire  _GEN_6769 = _T_49 ? _GEN_2092 : _GEN_6233; // @[dcache.scala 382:13]
  wire  _GEN_6770 = _T_49 ? _GEN_2093 : _GEN_6234; // @[dcache.scala 382:13]
  wire  _GEN_6771 = _T_49 ? _GEN_2094 : _GEN_6235; // @[dcache.scala 382:13]
  wire  _GEN_6772 = _T_49 ? _GEN_2095 : _GEN_6236; // @[dcache.scala 382:13]
  wire  _GEN_6773 = _T_49 ? _GEN_2096 : _GEN_6237; // @[dcache.scala 382:13]
  wire  _GEN_6774 = _T_49 ? _GEN_2097 : _GEN_6238; // @[dcache.scala 382:13]
  wire  _GEN_6775 = _T_49 ? _GEN_2098 : _GEN_6239; // @[dcache.scala 382:13]
  wire  _GEN_6776 = _T_49 ? _GEN_2099 : _GEN_6240; // @[dcache.scala 382:13]
  wire  _GEN_6777 = _T_49 ? _GEN_2100 : _GEN_6241; // @[dcache.scala 382:13]
  wire  _GEN_6778 = _T_49 ? _GEN_2101 : _GEN_6242; // @[dcache.scala 382:13]
  wire  _GEN_6779 = _T_49 ? _GEN_2102 : _GEN_6243; // @[dcache.scala 382:13]
  wire  _GEN_6780 = _T_49 ? _GEN_2103 : _GEN_6244; // @[dcache.scala 382:13]
  wire  _GEN_6781 = _T_49 ? _GEN_2104 : _GEN_6245; // @[dcache.scala 382:13]
  wire  _GEN_6782 = _T_49 ? _GEN_2105 : _GEN_6246; // @[dcache.scala 382:13]
  wire  _GEN_6783 = _T_49 ? _GEN_2106 : _GEN_6247; // @[dcache.scala 382:13]
  wire  _GEN_6784 = _T_49 ? _GEN_2107 : _GEN_6248; // @[dcache.scala 382:13]
  wire  _GEN_6785 = _T_49 ? _GEN_2108 : _GEN_6249; // @[dcache.scala 382:13]
  wire  _GEN_6786 = _T_49 ? _GEN_2109 : _GEN_6250; // @[dcache.scala 382:13]
  wire  _GEN_6787 = _T_49 ? _GEN_2110 : _GEN_6251; // @[dcache.scala 382:13]
  wire  _GEN_6788 = _T_49 ? _GEN_2111 : _GEN_6252; // @[dcache.scala 382:13]
  wire  _GEN_6789 = _T_49 ? _GEN_2112 : _GEN_6253; // @[dcache.scala 382:13]
  wire  _GEN_6790 = _T_49 ? _GEN_2113 : _GEN_6254; // @[dcache.scala 382:13]
  wire  _GEN_6791 = _T_49 ? _GEN_2114 : _GEN_6255; // @[dcache.scala 382:13]
  wire  _GEN_6792 = _T_49 ? _GEN_2115 : _GEN_6256; // @[dcache.scala 382:13]
  wire  _GEN_6793 = _T_49 ? _GEN_2116 : _GEN_6257; // @[dcache.scala 382:13]
  wire  _GEN_6794 = _T_49 ? _GEN_2117 : _GEN_6258; // @[dcache.scala 382:13]
  wire  _GEN_6795 = _T_49 ? _GEN_2118 : _GEN_6259; // @[dcache.scala 382:13]
  wire  _GEN_6796 = _T_49 ? _GEN_2119 : _GEN_6260; // @[dcache.scala 382:13]
  wire  _GEN_6797 = _T_49 ? _GEN_2120 : _GEN_6261; // @[dcache.scala 382:13]
  wire  _GEN_6798 = _T_49 ? _GEN_2121 : _GEN_6262; // @[dcache.scala 382:13]
  wire  _GEN_6799 = _T_49 ? _GEN_2122 : _GEN_6263; // @[dcache.scala 382:13]
  wire  _GEN_6800 = _T_49 ? _GEN_2123 : _GEN_6264; // @[dcache.scala 382:13]
  wire  _GEN_6801 = _T_49 ? _GEN_2124 : _GEN_6265; // @[dcache.scala 382:13]
  wire  _GEN_6802 = _T_49 ? _GEN_2125 : _GEN_6266; // @[dcache.scala 382:13]
  wire  _GEN_6803 = _T_49 ? _GEN_2126 : _GEN_6267; // @[dcache.scala 382:13]
  wire  _GEN_6804 = _T_49 ? _GEN_2127 : _GEN_6268; // @[dcache.scala 382:13]
  wire  _GEN_6805 = _T_49 ? _GEN_2128 : _GEN_6269; // @[dcache.scala 382:13]
  wire  _GEN_6806 = _T_49 ? _GEN_2129 : _GEN_6270; // @[dcache.scala 382:13]
  wire  _GEN_6807 = _T_49 ? _GEN_2130 : _GEN_6271; // @[dcache.scala 382:13]
  wire  _GEN_6808 = _T_49 ? _GEN_2131 : _GEN_6272; // @[dcache.scala 382:13]
  wire  _GEN_6809 = _T_49 ? _GEN_2132 : _GEN_6273; // @[dcache.scala 382:13]
  wire  _GEN_6810 = _T_49 ? _GEN_2133 : _GEN_6274; // @[dcache.scala 382:13]
  wire  _GEN_6811 = _T_49 ? _GEN_2134 : _GEN_6275; // @[dcache.scala 382:13]
  wire  _GEN_6812 = _T_49 ? _GEN_2135 : _GEN_6276; // @[dcache.scala 382:13]
  wire  _GEN_6813 = _T_49 ? _GEN_2136 : _GEN_6277; // @[dcache.scala 382:13]
  wire  _GEN_6814 = _T_49 ? _GEN_2137 : _GEN_6278; // @[dcache.scala 382:13]
  wire  _GEN_6815 = _T_49 ? _GEN_2138 : _GEN_6279; // @[dcache.scala 382:13]
  wire  _GEN_6816 = _T_49 ? _GEN_2139 : _GEN_6280; // @[dcache.scala 382:13]
  wire  _GEN_6817 = _T_49 ? _GEN_2140 : _GEN_6281; // @[dcache.scala 382:13]
  wire  _GEN_6818 = _T_49 ? _GEN_2141 : _GEN_6282; // @[dcache.scala 382:13]
  wire  _GEN_6819 = _T_49 ? _GEN_2142 : _GEN_6283; // @[dcache.scala 382:13]
  wire  _GEN_6820 = _T_49 ? _GEN_2143 : _GEN_6284; // @[dcache.scala 382:13]
  wire  _GEN_6821 = _T_49 ? _GEN_2144 : _GEN_6285; // @[dcache.scala 382:13]
  wire  _GEN_6822 = _T_49 ? _GEN_2145 : _GEN_6286; // @[dcache.scala 382:13]
  wire  _GEN_6823 = _T_49 ? _GEN_2146 : _GEN_6287; // @[dcache.scala 382:13]
  wire  _GEN_6824 = _T_49 ? _GEN_2147 : _GEN_6288; // @[dcache.scala 382:13]
  wire  _GEN_6825 = _T_49 ? _GEN_2148 : _GEN_6289; // @[dcache.scala 382:13]
  wire  _GEN_6826 = _T_49 ? _GEN_2149 : _GEN_6290; // @[dcache.scala 382:13]
  wire  _GEN_6827 = _T_49 ? _GEN_2150 : _GEN_6291; // @[dcache.scala 382:13]
  wire  _GEN_6828 = _T_49 ? _GEN_2151 : _GEN_6292; // @[dcache.scala 382:13]
  wire  _GEN_6829 = _T_49 ? _GEN_2152 : _GEN_6293; // @[dcache.scala 382:13]
  wire  _GEN_6830 = _T_49 ? _GEN_2153 : _GEN_6294; // @[dcache.scala 382:13]
  wire  _GEN_6831 = _T_49 ? _GEN_2154 : _GEN_6295; // @[dcache.scala 382:13]
  wire  _GEN_6832 = _T_49 ? _GEN_2155 : _GEN_6296; // @[dcache.scala 382:13]
  wire  _GEN_6833 = _T_49 ? _GEN_2156 : _GEN_6297; // @[dcache.scala 382:13]
  wire  _GEN_6834 = _T_49 ? _GEN_2157 : _GEN_6298; // @[dcache.scala 382:13]
  wire  _GEN_6835 = _T_49 ? _GEN_2158 : _GEN_6299; // @[dcache.scala 382:13]
  wire  _GEN_6836 = _T_49 ? _GEN_2159 : _GEN_6300; // @[dcache.scala 382:13]
  wire  _GEN_6837 = _T_49 ? _GEN_2160 : _GEN_6301; // @[dcache.scala 382:13]
  wire  _GEN_6838 = _T_49 ? _GEN_2161 : _GEN_6302; // @[dcache.scala 382:13]
  wire  _GEN_6839 = _T_49 ? _GEN_2162 : _GEN_6303; // @[dcache.scala 382:13]
  wire  _GEN_6840 = _T_49 ? _GEN_2163 : _GEN_6304; // @[dcache.scala 382:13]
  wire  _GEN_6841 = _T_49 ? _GEN_2164 : _GEN_6305; // @[dcache.scala 382:13]
  wire  _GEN_6842 = _T_49 ? _GEN_2165 : _GEN_6306; // @[dcache.scala 382:13]
  wire  _GEN_6843 = _T_49 ? _GEN_2166 : _GEN_6307; // @[dcache.scala 382:13]
  wire  _GEN_6844 = _T_49 ? _GEN_2167 : _GEN_6308; // @[dcache.scala 382:13]
  wire  _GEN_6845 = _T_49 ? _GEN_2168 : _GEN_6309; // @[dcache.scala 382:13]
  wire  _GEN_6846 = _T_49 ? _GEN_2169 : _GEN_6310; // @[dcache.scala 382:13]
  wire  _GEN_6847 = _T_49 ? _GEN_2170 : _GEN_6311; // @[dcache.scala 382:13]
  wire  _GEN_6848 = _T_49 ? _GEN_2171 : _GEN_6312; // @[dcache.scala 382:13]
  wire  _GEN_6849 = _T_49 ? _GEN_2172 : _GEN_6313; // @[dcache.scala 382:13]
  wire  _GEN_6850 = _T_49 ? _GEN_2173 : _GEN_6314; // @[dcache.scala 382:13]
  wire  _GEN_6851 = _T_49 ? _GEN_2174 : _GEN_6315; // @[dcache.scala 382:13]
  wire  _GEN_6852 = _T_49 ? _GEN_2175 : _GEN_6316; // @[dcache.scala 382:13]
  wire  _GEN_6853 = _T_49 ? _GEN_2176 : _GEN_6317; // @[dcache.scala 382:13]
  wire  _GEN_6854 = _T_49 ? _GEN_2177 : _GEN_6318; // @[dcache.scala 382:13]
  wire  _GEN_6855 = _T_49 ? _GEN_2178 : _GEN_6319; // @[dcache.scala 382:13]
  wire  _GEN_6856 = _T_49 ? _GEN_2179 : _GEN_6320; // @[dcache.scala 382:13]
  wire  _GEN_6857 = _T_49 ? _GEN_2180 : _GEN_6321; // @[dcache.scala 382:13]
  wire  _GEN_6858 = _T_49 ? _GEN_2181 : _GEN_6322; // @[dcache.scala 382:13]
  wire  _GEN_6859 = _T_49 ? _GEN_2182 : _GEN_6323; // @[dcache.scala 382:13]
  wire  _GEN_6860 = _T_49 ? _GEN_2183 : _GEN_6324; // @[dcache.scala 382:13]
  wire  _GEN_6861 = _T_49 ? _GEN_2184 : _GEN_6325; // @[dcache.scala 382:13]
  wire  _GEN_6862 = _T_49 ? _GEN_2185 : _GEN_6326; // @[dcache.scala 382:13]
  wire  _GEN_6863 = _T_49 ? _GEN_2186 : _GEN_6327; // @[dcache.scala 382:13]
  wire  _GEN_6864 = _T_49 ? _GEN_2187 : _GEN_6328; // @[dcache.scala 382:13]
  wire  _GEN_6865 = _T_49 ? _GEN_2188 : _GEN_6329; // @[dcache.scala 382:13]
  wire  _GEN_6866 = _T_49 ? _GEN_2189 : _GEN_6330; // @[dcache.scala 382:13]
  wire  _GEN_6867 = _T_49 ? _GEN_2190 : _GEN_6331; // @[dcache.scala 382:13]
  wire  _GEN_6868 = _T_49 ? _GEN_2191 : _GEN_6332; // @[dcache.scala 382:13]
  wire  _GEN_6869 = _T_49 ? _GEN_2192 : _GEN_6333; // @[dcache.scala 382:13]
  wire  _GEN_6870 = _T_49 ? _GEN_2193 : _GEN_6334; // @[dcache.scala 382:13]
  wire  _GEN_6871 = _T_49 ? _GEN_2194 : _GEN_6335; // @[dcache.scala 382:13]
  wire  _GEN_6872 = _T_49 ? _GEN_2195 : _GEN_6336; // @[dcache.scala 382:13]
  wire  _GEN_6873 = _T_49 ? _GEN_2196 : _GEN_6337; // @[dcache.scala 382:13]
  wire  _GEN_6874 = _T_49 ? _GEN_2197 : _GEN_6338; // @[dcache.scala 382:13]
  wire  _GEN_6875 = _T_49 ? _GEN_2198 : _GEN_6339; // @[dcache.scala 382:13]
  wire  _GEN_6876 = _T_49 ? _GEN_2199 : _GEN_6340; // @[dcache.scala 382:13]
  wire  _GEN_6877 = _T_49 ? _GEN_2200 : _GEN_6341; // @[dcache.scala 382:13]
  wire  _GEN_6878 = _T_49 ? _GEN_2201 : _GEN_6342; // @[dcache.scala 382:13]
  wire  _GEN_6879 = _T_49 ? _GEN_2202 : _GEN_6343; // @[dcache.scala 382:13]
  wire  _GEN_6880 = _T_49 ? _GEN_2203 : _GEN_6344; // @[dcache.scala 382:13]
  wire  _GEN_6881 = _T_49 ? _GEN_2204 : _GEN_6345; // @[dcache.scala 382:13]
  wire  _GEN_6882 = _T_49 ? _GEN_2205 : _GEN_6346; // @[dcache.scala 382:13]
  wire  _GEN_6883 = _T_49 ? _GEN_2206 : _GEN_6347; // @[dcache.scala 382:13]
  wire  _GEN_6884 = _T_49 ? _GEN_2207 : _GEN_6348; // @[dcache.scala 382:13]
  wire  _GEN_6885 = _T_49 ? _GEN_2208 : _GEN_6349; // @[dcache.scala 382:13]
  wire  _GEN_6886 = _T_49 ? _GEN_2209 : _GEN_6350; // @[dcache.scala 382:13]
  wire  _GEN_6887 = _T_49 ? _GEN_2210 : _GEN_6351; // @[dcache.scala 382:13]
  wire  _GEN_6888 = _T_49 ? _GEN_2211 : _GEN_6352; // @[dcache.scala 382:13]
  wire  _GEN_6889 = _T_49 ? _GEN_2212 : _GEN_6353; // @[dcache.scala 382:13]
  wire  _GEN_6890 = _T_49 ? _GEN_2213 : _GEN_6354; // @[dcache.scala 382:13]
  wire  _GEN_6891 = _T_49 ? _GEN_2214 : _GEN_6355; // @[dcache.scala 382:13]
  wire  _GEN_6892 = _T_49 ? _GEN_2215 : _GEN_6356; // @[dcache.scala 382:13]
  wire  _GEN_6893 = _T_49 ? _GEN_2216 : _GEN_6357; // @[dcache.scala 382:13]
  wire  _GEN_6894 = _T_49 ? _GEN_2217 : _GEN_6358; // @[dcache.scala 382:13]
  wire  _GEN_6895 = _T_49 ? _GEN_2218 : _GEN_6359; // @[dcache.scala 382:13]
  wire  _GEN_6896 = _T_49 ? _GEN_2219 : _GEN_6360; // @[dcache.scala 382:13]
  wire  _GEN_6897 = _T_49 ? _GEN_2220 : _GEN_6361; // @[dcache.scala 382:13]
  wire  _GEN_6898 = _T_49 ? _GEN_2221 : _GEN_6362; // @[dcache.scala 382:13]
  wire  _GEN_6899 = _T_49 ? _GEN_2222 : _GEN_6363; // @[dcache.scala 382:13]
  wire  _GEN_6900 = _T_49 ? _GEN_2223 : _GEN_6364; // @[dcache.scala 382:13]
  wire  _GEN_6901 = _T_49 ? _GEN_2224 : _GEN_6365; // @[dcache.scala 382:13]
  wire  _GEN_6902 = _T_49 ? _GEN_2225 : _GEN_6366; // @[dcache.scala 382:13]
  wire  _GEN_6903 = _T_49 ? _GEN_2226 : _GEN_6367; // @[dcache.scala 382:13]
  wire  _GEN_6904 = _T_49 ? _GEN_2227 : _GEN_6368; // @[dcache.scala 382:13]
  wire  _GEN_6905 = _T_49 ? _GEN_2228 : _GEN_6369; // @[dcache.scala 382:13]
  wire  _GEN_6906 = _T_49 ? _GEN_2229 : _GEN_6370; // @[dcache.scala 382:13]
  wire  _GEN_6907 = _T_49 ? _GEN_2230 : _GEN_6371; // @[dcache.scala 382:13]
  wire  _GEN_6908 = _T_49 ? _GEN_2231 : _GEN_6372; // @[dcache.scala 382:13]
  wire  _GEN_6909 = _T_49 ? _GEN_2232 : _GEN_6373; // @[dcache.scala 382:13]
  wire  _GEN_6910 = _T_49 ? _GEN_2233 : _GEN_6374; // @[dcache.scala 382:13]
  wire  _GEN_6911 = _T_49 ? _GEN_2234 : _GEN_6375; // @[dcache.scala 382:13]
  wire  _GEN_6912 = _T_49 ? _GEN_2235 : _GEN_6376; // @[dcache.scala 382:13]
  wire  _GEN_6913 = _T_49 ? _GEN_2236 : _GEN_6377; // @[dcache.scala 382:13]
  wire  _GEN_6914 = _T_49 ? _GEN_2237 : _GEN_6378; // @[dcache.scala 382:13]
  wire  _GEN_6915 = _T_49 ? _GEN_2238 : _GEN_6379; // @[dcache.scala 382:13]
  wire  _GEN_6916 = _T_49 ? _GEN_2239 : _GEN_6380; // @[dcache.scala 382:13]
  wire  _GEN_6917 = _T_49 ? _GEN_2240 : _GEN_6381; // @[dcache.scala 382:13]
  wire  _GEN_6918 = _T_49 ? _GEN_2241 : _GEN_6382; // @[dcache.scala 382:13]
  wire  _GEN_6919 = _T_49 ? _GEN_2242 : _GEN_6383; // @[dcache.scala 382:13]
  wire  _GEN_6920 = _T_49 ? _GEN_2243 : _GEN_6384; // @[dcache.scala 382:13]
  wire  _GEN_6921 = _T_49 ? _GEN_2244 : _GEN_6385; // @[dcache.scala 382:13]
  wire  _GEN_6922 = _T_49 ? _GEN_2245 : _GEN_6386; // @[dcache.scala 382:13]
  wire  _GEN_6923 = _T_49 ? _GEN_2246 : _GEN_6387; // @[dcache.scala 382:13]
  wire  _GEN_6924 = _T_49 ? _GEN_2247 : _GEN_6388; // @[dcache.scala 382:13]
  wire  _GEN_6925 = _T_49 ? _GEN_2248 : _GEN_6389; // @[dcache.scala 382:13]
  wire  _GEN_6926 = _T_49 ? _GEN_2249 : _GEN_6390; // @[dcache.scala 382:13]
  wire  _GEN_6927 = _T_49 ? _GEN_2250 : _GEN_6391; // @[dcache.scala 382:13]
  wire  _GEN_6928 = _T_49 ? _GEN_2251 : _GEN_6392; // @[dcache.scala 382:13]
  wire  _GEN_6929 = _T_49 ? _GEN_2252 : _GEN_6393; // @[dcache.scala 382:13]
  wire  _GEN_6930 = _T_49 ? _GEN_2253 : _GEN_6394; // @[dcache.scala 382:13]
  wire  _GEN_6931 = _T_49 ? _GEN_2254 : _GEN_6395; // @[dcache.scala 382:13]
  wire  _GEN_6932 = _T_49 ? _GEN_2255 : _GEN_6396; // @[dcache.scala 382:13]
  wire  _GEN_6933 = _T_49 ? _GEN_2256 : _GEN_6397; // @[dcache.scala 382:13]
  wire  _GEN_6934 = _T_49 ? _GEN_2257 : _GEN_6398; // @[dcache.scala 382:13]
  wire  _GEN_6935 = _T_49 ? _GEN_2258 : _GEN_6399; // @[dcache.scala 382:13]
  wire  _GEN_6936 = _T_49 ? _GEN_2259 : _GEN_6400; // @[dcache.scala 382:13]
  wire  _GEN_6937 = _T_49 ? _GEN_2260 : _GEN_6401; // @[dcache.scala 382:13]
  wire  _GEN_6938 = _T_49 ? _GEN_2261 : _GEN_6402; // @[dcache.scala 382:13]
  wire  _GEN_6939 = _T_49 ? _GEN_2262 : _GEN_6403; // @[dcache.scala 382:13]
  wire  _GEN_6940 = _T_49 ? _GEN_2263 : _GEN_6404; // @[dcache.scala 382:13]
  wire  _GEN_6941 = _T_49 ? _GEN_2264 : _GEN_6405; // @[dcache.scala 382:13]
  wire  _GEN_6942 = _T_49 ? _GEN_2265 : _GEN_6406; // @[dcache.scala 382:13]
  wire  _GEN_6943 = _T_49 ? _GEN_2266 : _GEN_6407; // @[dcache.scala 382:13]
  wire  _GEN_6944 = _T_49 ? _GEN_2267 : _GEN_6408; // @[dcache.scala 382:13]
  wire  _GEN_6945 = _T_49 ? _GEN_2268 : _GEN_6409; // @[dcache.scala 382:13]
  wire  _GEN_6946 = _T_49 ? _GEN_2269 : _GEN_6410; // @[dcache.scala 382:13]
  wire  _GEN_6947 = _T_49 ? _GEN_2270 : _GEN_6411; // @[dcache.scala 382:13]
  wire  _GEN_6948 = _T_49 ? _GEN_2271 : _GEN_6412; // @[dcache.scala 382:13]
  wire  _GEN_6949 = _T_49 ? _GEN_2272 : _GEN_6413; // @[dcache.scala 382:13]
  wire  _GEN_6950 = _T_49 ? _GEN_2273 : _GEN_6414; // @[dcache.scala 382:13]
  wire  _GEN_6951 = _T_49 ? _GEN_2274 : _GEN_6415; // @[dcache.scala 382:13]
  wire  _GEN_6952 = _T_49 ? _GEN_2275 : _GEN_6416; // @[dcache.scala 382:13]
  wire  _GEN_6953 = _T_49 ? _GEN_2276 : _GEN_6417; // @[dcache.scala 382:13]
  wire  _GEN_6954 = _T_49 ? _GEN_2277 : _GEN_6418; // @[dcache.scala 382:13]
  wire  _GEN_6955 = _T_49 ? _GEN_2278 : _GEN_6419; // @[dcache.scala 382:13]
  wire  _GEN_6956 = _T_49 ? _GEN_2279 : _GEN_6420; // @[dcache.scala 382:13]
  wire  _GEN_6957 = _T_49 ? _GEN_2280 : _GEN_6421; // @[dcache.scala 382:13]
  wire  _GEN_6958 = _T_49 ? _GEN_2281 : _GEN_6422; // @[dcache.scala 382:13]
  wire  _GEN_6959 = _T_49 ? _GEN_2282 : _GEN_6423; // @[dcache.scala 382:13]
  wire  _GEN_6960 = _T_49 ? _GEN_2283 : _GEN_6424; // @[dcache.scala 382:13]
  wire  _GEN_6961 = _T_49 ? _GEN_2284 : _GEN_6425; // @[dcache.scala 382:13]
  wire  _GEN_6962 = _T_49 ? _GEN_2285 : _GEN_6426; // @[dcache.scala 382:13]
  wire  _GEN_6963 = _T_49 ? _GEN_2286 : _GEN_6427; // @[dcache.scala 382:13]
  wire  _GEN_6964 = _T_49 ? _GEN_2287 : _GEN_6428; // @[dcache.scala 382:13]
  wire  _GEN_6965 = _T_49 ? _GEN_2288 : _GEN_6429; // @[dcache.scala 382:13]
  wire  _GEN_6966 = _T_49 ? _GEN_2289 : _GEN_6430; // @[dcache.scala 382:13]
  wire  _GEN_6967 = _T_49 ? _GEN_2290 : _GEN_6431; // @[dcache.scala 382:13]
  wire  _GEN_6968 = _T_49 ? _GEN_2291 : _GEN_6432; // @[dcache.scala 382:13]
  wire  _GEN_6969 = _T_49 ? _GEN_2292 : _GEN_6433; // @[dcache.scala 382:13]
  wire  _GEN_6970 = _T_49 ? _GEN_2293 : _GEN_6434; // @[dcache.scala 382:13]
  wire  _GEN_6971 = _T_49 ? _GEN_2294 : _GEN_6435; // @[dcache.scala 382:13]
  wire  _GEN_6972 = _T_49 ? _GEN_2295 : _GEN_6436; // @[dcache.scala 382:13]
  wire  _GEN_6973 = _T_49 ? _GEN_2296 : _GEN_5923; // @[dcache.scala 382:13]
  wire  _GEN_6974 = _T_49 ? _GEN_2297 : _GEN_5924; // @[dcache.scala 382:13]
  wire [20:0] _GEN_6975 = _T_49 ? _GEN_2298 : _GEN_5921; // @[dcache.scala 382:13]
  wire [20:0] _GEN_6976 = _T_49 ? _GEN_2299 : _GEN_5922; // @[dcache.scala 382:13]
  wire  _GEN_6977 = _T_49 ? 1'h0 : _GEN_5915; // @[dcache.scala 382:13 157:25]
  wire [31:0] _GEN_6978 = _T_49 ? 32'h7777 : _GEN_5916; // @[dcache.scala 382:13 155:25]
  wire  _GEN_6979 = _T_49 ? req_valid : _GEN_5918; // @[dcache.scala 382:13 116:34]
  wire  _GEN_6980 = _T_49 ? 1'h0 : _GEN_5919; // @[dcache.scala 382:13 97:21]
  wire [21:0] _GEN_6981 = _T_49 ? 22'h0 : _GEN_5920; // @[dcache.scala 382:13 98:21]
  wire  _GEN_6982 = _T_49 ? cacheInst_r : _GEN_6437; // @[dcache.scala 382:13 89:38]
  wire  _GEN_6983 = _T_49 ? invalidate : _GEN_6438; // @[dcache.scala 382:13 90:38]
  wire  _GEN_6984 = _T_49 ? indexOnly : _GEN_6439; // @[dcache.scala 382:13 94:38]
  wire  _GEN_6985 = _T_49 ? writeBack : _GEN_6440; // @[dcache.scala 382:13 93:38]
  wire  _GEN_6986 = _T_49 ? storeTag : _GEN_6441; // @[dcache.scala 382:13 92:38]
  wire  _GEN_6987 = _T_49 ? loadTag : _GEN_6442; // @[dcache.scala 382:13 91:38]
  wire [2:0] _GEN_6988 = 3'h5 == state ? _GEN_6460 : state; // @[dcache.scala 183:18 171:34]
  wire [1:0] _GEN_6989 = 3'h5 == state ? _GEN_6443 : wr_cnt; // @[dcache.scala 183:18 178:34]
  wire [31:0] _GEN_6990 = 3'h5 == state ? _GEN_6444 : 32'h0; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_6991 = 3'h5 == state ? _GEN_6445 : 32'h0; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_6992 = 3'h5 == state ? _GEN_6446 : 32'h0; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_6993 = 3'h5 == state ? _GEN_6447 : 32'h0; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_6994 = 3'h5 == state ? _GEN_6448 : 32'h0; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_6995 = 3'h5 == state ? _GEN_6449 : 32'h0; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_6996 = 3'h5 == state ? _GEN_6450 : 32'h0; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_6997 = 3'h5 == state ? _GEN_6451 : 32'h0; // @[dcache.scala 183:18 149:33]
  wire [3:0] _GEN_6998 = 3'h5 == state ? _GEN_6452 : 4'h0; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_6999 = 3'h5 == state ? _GEN_6453 : 4'h0; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7000 = 3'h5 == state ? _GEN_6454 : 4'h0; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7001 = 3'h5 == state ? _GEN_6455 : 4'h0; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7002 = 3'h5 == state ? _GEN_6456 : 4'h0; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7003 = 3'h5 == state ? _GEN_6457 : 4'h0; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7004 = 3'h5 == state ? _GEN_6458 : 4'h0; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7005 = 3'h5 == state ? _GEN_6459 : 4'h0; // @[dcache.scala 183:18 150:33]
  wire  _GEN_7006 = 3'h5 == state ? _GEN_6461 : dirty_0_0; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7007 = 3'h5 == state ? _GEN_6462 : dirty_0_1; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7008 = 3'h5 == state ? _GEN_6463 : dirty_0_2; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7009 = 3'h5 == state ? _GEN_6464 : dirty_0_3; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7010 = 3'h5 == state ? _GEN_6465 : dirty_0_4; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7011 = 3'h5 == state ? _GEN_6466 : dirty_0_5; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7012 = 3'h5 == state ? _GEN_6467 : dirty_0_6; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7013 = 3'h5 == state ? _GEN_6468 : dirty_0_7; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7014 = 3'h5 == state ? _GEN_6469 : dirty_0_8; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7015 = 3'h5 == state ? _GEN_6470 : dirty_0_9; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7016 = 3'h5 == state ? _GEN_6471 : dirty_0_10; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7017 = 3'h5 == state ? _GEN_6472 : dirty_0_11; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7018 = 3'h5 == state ? _GEN_6473 : dirty_0_12; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7019 = 3'h5 == state ? _GEN_6474 : dirty_0_13; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7020 = 3'h5 == state ? _GEN_6475 : dirty_0_14; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7021 = 3'h5 == state ? _GEN_6476 : dirty_0_15; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7022 = 3'h5 == state ? _GEN_6477 : dirty_0_16; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7023 = 3'h5 == state ? _GEN_6478 : dirty_0_17; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7024 = 3'h5 == state ? _GEN_6479 : dirty_0_18; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7025 = 3'h5 == state ? _GEN_6480 : dirty_0_19; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7026 = 3'h5 == state ? _GEN_6481 : dirty_0_20; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7027 = 3'h5 == state ? _GEN_6482 : dirty_0_21; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7028 = 3'h5 == state ? _GEN_6483 : dirty_0_22; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7029 = 3'h5 == state ? _GEN_6484 : dirty_0_23; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7030 = 3'h5 == state ? _GEN_6485 : dirty_0_24; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7031 = 3'h5 == state ? _GEN_6486 : dirty_0_25; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7032 = 3'h5 == state ? _GEN_6487 : dirty_0_26; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7033 = 3'h5 == state ? _GEN_6488 : dirty_0_27; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7034 = 3'h5 == state ? _GEN_6489 : dirty_0_28; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7035 = 3'h5 == state ? _GEN_6490 : dirty_0_29; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7036 = 3'h5 == state ? _GEN_6491 : dirty_0_30; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7037 = 3'h5 == state ? _GEN_6492 : dirty_0_31; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7038 = 3'h5 == state ? _GEN_6493 : dirty_0_32; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7039 = 3'h5 == state ? _GEN_6494 : dirty_0_33; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7040 = 3'h5 == state ? _GEN_6495 : dirty_0_34; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7041 = 3'h5 == state ? _GEN_6496 : dirty_0_35; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7042 = 3'h5 == state ? _GEN_6497 : dirty_0_36; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7043 = 3'h5 == state ? _GEN_6498 : dirty_0_37; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7044 = 3'h5 == state ? _GEN_6499 : dirty_0_38; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7045 = 3'h5 == state ? _GEN_6500 : dirty_0_39; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7046 = 3'h5 == state ? _GEN_6501 : dirty_0_40; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7047 = 3'h5 == state ? _GEN_6502 : dirty_0_41; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7048 = 3'h5 == state ? _GEN_6503 : dirty_0_42; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7049 = 3'h5 == state ? _GEN_6504 : dirty_0_43; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7050 = 3'h5 == state ? _GEN_6505 : dirty_0_44; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7051 = 3'h5 == state ? _GEN_6506 : dirty_0_45; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7052 = 3'h5 == state ? _GEN_6507 : dirty_0_46; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7053 = 3'h5 == state ? _GEN_6508 : dirty_0_47; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7054 = 3'h5 == state ? _GEN_6509 : dirty_0_48; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7055 = 3'h5 == state ? _GEN_6510 : dirty_0_49; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7056 = 3'h5 == state ? _GEN_6511 : dirty_0_50; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7057 = 3'h5 == state ? _GEN_6512 : dirty_0_51; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7058 = 3'h5 == state ? _GEN_6513 : dirty_0_52; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7059 = 3'h5 == state ? _GEN_6514 : dirty_0_53; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7060 = 3'h5 == state ? _GEN_6515 : dirty_0_54; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7061 = 3'h5 == state ? _GEN_6516 : dirty_0_55; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7062 = 3'h5 == state ? _GEN_6517 : dirty_0_56; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7063 = 3'h5 == state ? _GEN_6518 : dirty_0_57; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7064 = 3'h5 == state ? _GEN_6519 : dirty_0_58; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7065 = 3'h5 == state ? _GEN_6520 : dirty_0_59; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7066 = 3'h5 == state ? _GEN_6521 : dirty_0_60; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7067 = 3'h5 == state ? _GEN_6522 : dirty_0_61; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7068 = 3'h5 == state ? _GEN_6523 : dirty_0_62; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7069 = 3'h5 == state ? _GEN_6524 : dirty_0_63; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7070 = 3'h5 == state ? _GEN_6525 : dirty_0_64; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7071 = 3'h5 == state ? _GEN_6526 : dirty_0_65; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7072 = 3'h5 == state ? _GEN_6527 : dirty_0_66; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7073 = 3'h5 == state ? _GEN_6528 : dirty_0_67; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7074 = 3'h5 == state ? _GEN_6529 : dirty_0_68; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7075 = 3'h5 == state ? _GEN_6530 : dirty_0_69; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7076 = 3'h5 == state ? _GEN_6531 : dirty_0_70; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7077 = 3'h5 == state ? _GEN_6532 : dirty_0_71; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7078 = 3'h5 == state ? _GEN_6533 : dirty_0_72; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7079 = 3'h5 == state ? _GEN_6534 : dirty_0_73; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7080 = 3'h5 == state ? _GEN_6535 : dirty_0_74; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7081 = 3'h5 == state ? _GEN_6536 : dirty_0_75; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7082 = 3'h5 == state ? _GEN_6537 : dirty_0_76; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7083 = 3'h5 == state ? _GEN_6538 : dirty_0_77; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7084 = 3'h5 == state ? _GEN_6539 : dirty_0_78; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7085 = 3'h5 == state ? _GEN_6540 : dirty_0_79; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7086 = 3'h5 == state ? _GEN_6541 : dirty_0_80; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7087 = 3'h5 == state ? _GEN_6542 : dirty_0_81; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7088 = 3'h5 == state ? _GEN_6543 : dirty_0_82; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7089 = 3'h5 == state ? _GEN_6544 : dirty_0_83; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7090 = 3'h5 == state ? _GEN_6545 : dirty_0_84; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7091 = 3'h5 == state ? _GEN_6546 : dirty_0_85; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7092 = 3'h5 == state ? _GEN_6547 : dirty_0_86; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7093 = 3'h5 == state ? _GEN_6548 : dirty_0_87; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7094 = 3'h5 == state ? _GEN_6549 : dirty_0_88; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7095 = 3'h5 == state ? _GEN_6550 : dirty_0_89; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7096 = 3'h5 == state ? _GEN_6551 : dirty_0_90; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7097 = 3'h5 == state ? _GEN_6552 : dirty_0_91; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7098 = 3'h5 == state ? _GEN_6553 : dirty_0_92; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7099 = 3'h5 == state ? _GEN_6554 : dirty_0_93; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7100 = 3'h5 == state ? _GEN_6555 : dirty_0_94; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7101 = 3'h5 == state ? _GEN_6556 : dirty_0_95; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7102 = 3'h5 == state ? _GEN_6557 : dirty_0_96; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7103 = 3'h5 == state ? _GEN_6558 : dirty_0_97; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7104 = 3'h5 == state ? _GEN_6559 : dirty_0_98; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7105 = 3'h5 == state ? _GEN_6560 : dirty_0_99; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7106 = 3'h5 == state ? _GEN_6561 : dirty_0_100; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7107 = 3'h5 == state ? _GEN_6562 : dirty_0_101; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7108 = 3'h5 == state ? _GEN_6563 : dirty_0_102; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7109 = 3'h5 == state ? _GEN_6564 : dirty_0_103; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7110 = 3'h5 == state ? _GEN_6565 : dirty_0_104; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7111 = 3'h5 == state ? _GEN_6566 : dirty_0_105; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7112 = 3'h5 == state ? _GEN_6567 : dirty_0_106; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7113 = 3'h5 == state ? _GEN_6568 : dirty_0_107; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7114 = 3'h5 == state ? _GEN_6569 : dirty_0_108; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7115 = 3'h5 == state ? _GEN_6570 : dirty_0_109; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7116 = 3'h5 == state ? _GEN_6571 : dirty_0_110; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7117 = 3'h5 == state ? _GEN_6572 : dirty_0_111; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7118 = 3'h5 == state ? _GEN_6573 : dirty_0_112; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7119 = 3'h5 == state ? _GEN_6574 : dirty_0_113; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7120 = 3'h5 == state ? _GEN_6575 : dirty_0_114; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7121 = 3'h5 == state ? _GEN_6576 : dirty_0_115; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7122 = 3'h5 == state ? _GEN_6577 : dirty_0_116; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7123 = 3'h5 == state ? _GEN_6578 : dirty_0_117; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7124 = 3'h5 == state ? _GEN_6579 : dirty_0_118; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7125 = 3'h5 == state ? _GEN_6580 : dirty_0_119; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7126 = 3'h5 == state ? _GEN_6581 : dirty_0_120; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7127 = 3'h5 == state ? _GEN_6582 : dirty_0_121; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7128 = 3'h5 == state ? _GEN_6583 : dirty_0_122; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7129 = 3'h5 == state ? _GEN_6584 : dirty_0_123; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7130 = 3'h5 == state ? _GEN_6585 : dirty_0_124; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7131 = 3'h5 == state ? _GEN_6586 : dirty_0_125; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7132 = 3'h5 == state ? _GEN_6587 : dirty_0_126; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7133 = 3'h5 == state ? _GEN_6588 : dirty_0_127; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7134 = 3'h5 == state ? _GEN_6589 : dirty_0_128; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7135 = 3'h5 == state ? _GEN_6590 : dirty_0_129; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7136 = 3'h5 == state ? _GEN_6591 : dirty_0_130; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7137 = 3'h5 == state ? _GEN_6592 : dirty_0_131; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7138 = 3'h5 == state ? _GEN_6593 : dirty_0_132; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7139 = 3'h5 == state ? _GEN_6594 : dirty_0_133; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7140 = 3'h5 == state ? _GEN_6595 : dirty_0_134; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7141 = 3'h5 == state ? _GEN_6596 : dirty_0_135; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7142 = 3'h5 == state ? _GEN_6597 : dirty_0_136; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7143 = 3'h5 == state ? _GEN_6598 : dirty_0_137; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7144 = 3'h5 == state ? _GEN_6599 : dirty_0_138; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7145 = 3'h5 == state ? _GEN_6600 : dirty_0_139; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7146 = 3'h5 == state ? _GEN_6601 : dirty_0_140; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7147 = 3'h5 == state ? _GEN_6602 : dirty_0_141; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7148 = 3'h5 == state ? _GEN_6603 : dirty_0_142; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7149 = 3'h5 == state ? _GEN_6604 : dirty_0_143; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7150 = 3'h5 == state ? _GEN_6605 : dirty_0_144; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7151 = 3'h5 == state ? _GEN_6606 : dirty_0_145; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7152 = 3'h5 == state ? _GEN_6607 : dirty_0_146; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7153 = 3'h5 == state ? _GEN_6608 : dirty_0_147; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7154 = 3'h5 == state ? _GEN_6609 : dirty_0_148; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7155 = 3'h5 == state ? _GEN_6610 : dirty_0_149; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7156 = 3'h5 == state ? _GEN_6611 : dirty_0_150; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7157 = 3'h5 == state ? _GEN_6612 : dirty_0_151; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7158 = 3'h5 == state ? _GEN_6613 : dirty_0_152; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7159 = 3'h5 == state ? _GEN_6614 : dirty_0_153; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7160 = 3'h5 == state ? _GEN_6615 : dirty_0_154; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7161 = 3'h5 == state ? _GEN_6616 : dirty_0_155; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7162 = 3'h5 == state ? _GEN_6617 : dirty_0_156; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7163 = 3'h5 == state ? _GEN_6618 : dirty_0_157; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7164 = 3'h5 == state ? _GEN_6619 : dirty_0_158; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7165 = 3'h5 == state ? _GEN_6620 : dirty_0_159; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7166 = 3'h5 == state ? _GEN_6621 : dirty_0_160; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7167 = 3'h5 == state ? _GEN_6622 : dirty_0_161; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7168 = 3'h5 == state ? _GEN_6623 : dirty_0_162; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7169 = 3'h5 == state ? _GEN_6624 : dirty_0_163; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7170 = 3'h5 == state ? _GEN_6625 : dirty_0_164; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7171 = 3'h5 == state ? _GEN_6626 : dirty_0_165; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7172 = 3'h5 == state ? _GEN_6627 : dirty_0_166; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7173 = 3'h5 == state ? _GEN_6628 : dirty_0_167; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7174 = 3'h5 == state ? _GEN_6629 : dirty_0_168; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7175 = 3'h5 == state ? _GEN_6630 : dirty_0_169; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7176 = 3'h5 == state ? _GEN_6631 : dirty_0_170; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7177 = 3'h5 == state ? _GEN_6632 : dirty_0_171; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7178 = 3'h5 == state ? _GEN_6633 : dirty_0_172; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7179 = 3'h5 == state ? _GEN_6634 : dirty_0_173; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7180 = 3'h5 == state ? _GEN_6635 : dirty_0_174; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7181 = 3'h5 == state ? _GEN_6636 : dirty_0_175; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7182 = 3'h5 == state ? _GEN_6637 : dirty_0_176; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7183 = 3'h5 == state ? _GEN_6638 : dirty_0_177; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7184 = 3'h5 == state ? _GEN_6639 : dirty_0_178; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7185 = 3'h5 == state ? _GEN_6640 : dirty_0_179; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7186 = 3'h5 == state ? _GEN_6641 : dirty_0_180; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7187 = 3'h5 == state ? _GEN_6642 : dirty_0_181; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7188 = 3'h5 == state ? _GEN_6643 : dirty_0_182; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7189 = 3'h5 == state ? _GEN_6644 : dirty_0_183; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7190 = 3'h5 == state ? _GEN_6645 : dirty_0_184; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7191 = 3'h5 == state ? _GEN_6646 : dirty_0_185; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7192 = 3'h5 == state ? _GEN_6647 : dirty_0_186; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7193 = 3'h5 == state ? _GEN_6648 : dirty_0_187; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7194 = 3'h5 == state ? _GEN_6649 : dirty_0_188; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7195 = 3'h5 == state ? _GEN_6650 : dirty_0_189; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7196 = 3'h5 == state ? _GEN_6651 : dirty_0_190; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7197 = 3'h5 == state ? _GEN_6652 : dirty_0_191; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7198 = 3'h5 == state ? _GEN_6653 : dirty_0_192; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7199 = 3'h5 == state ? _GEN_6654 : dirty_0_193; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7200 = 3'h5 == state ? _GEN_6655 : dirty_0_194; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7201 = 3'h5 == state ? _GEN_6656 : dirty_0_195; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7202 = 3'h5 == state ? _GEN_6657 : dirty_0_196; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7203 = 3'h5 == state ? _GEN_6658 : dirty_0_197; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7204 = 3'h5 == state ? _GEN_6659 : dirty_0_198; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7205 = 3'h5 == state ? _GEN_6660 : dirty_0_199; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7206 = 3'h5 == state ? _GEN_6661 : dirty_0_200; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7207 = 3'h5 == state ? _GEN_6662 : dirty_0_201; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7208 = 3'h5 == state ? _GEN_6663 : dirty_0_202; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7209 = 3'h5 == state ? _GEN_6664 : dirty_0_203; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7210 = 3'h5 == state ? _GEN_6665 : dirty_0_204; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7211 = 3'h5 == state ? _GEN_6666 : dirty_0_205; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7212 = 3'h5 == state ? _GEN_6667 : dirty_0_206; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7213 = 3'h5 == state ? _GEN_6668 : dirty_0_207; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7214 = 3'h5 == state ? _GEN_6669 : dirty_0_208; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7215 = 3'h5 == state ? _GEN_6670 : dirty_0_209; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7216 = 3'h5 == state ? _GEN_6671 : dirty_0_210; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7217 = 3'h5 == state ? _GEN_6672 : dirty_0_211; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7218 = 3'h5 == state ? _GEN_6673 : dirty_0_212; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7219 = 3'h5 == state ? _GEN_6674 : dirty_0_213; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7220 = 3'h5 == state ? _GEN_6675 : dirty_0_214; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7221 = 3'h5 == state ? _GEN_6676 : dirty_0_215; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7222 = 3'h5 == state ? _GEN_6677 : dirty_0_216; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7223 = 3'h5 == state ? _GEN_6678 : dirty_0_217; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7224 = 3'h5 == state ? _GEN_6679 : dirty_0_218; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7225 = 3'h5 == state ? _GEN_6680 : dirty_0_219; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7226 = 3'h5 == state ? _GEN_6681 : dirty_0_220; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7227 = 3'h5 == state ? _GEN_6682 : dirty_0_221; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7228 = 3'h5 == state ? _GEN_6683 : dirty_0_222; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7229 = 3'h5 == state ? _GEN_6684 : dirty_0_223; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7230 = 3'h5 == state ? _GEN_6685 : dirty_0_224; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7231 = 3'h5 == state ? _GEN_6686 : dirty_0_225; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7232 = 3'h5 == state ? _GEN_6687 : dirty_0_226; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7233 = 3'h5 == state ? _GEN_6688 : dirty_0_227; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7234 = 3'h5 == state ? _GEN_6689 : dirty_0_228; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7235 = 3'h5 == state ? _GEN_6690 : dirty_0_229; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7236 = 3'h5 == state ? _GEN_6691 : dirty_0_230; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7237 = 3'h5 == state ? _GEN_6692 : dirty_0_231; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7238 = 3'h5 == state ? _GEN_6693 : dirty_0_232; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7239 = 3'h5 == state ? _GEN_6694 : dirty_0_233; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7240 = 3'h5 == state ? _GEN_6695 : dirty_0_234; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7241 = 3'h5 == state ? _GEN_6696 : dirty_0_235; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7242 = 3'h5 == state ? _GEN_6697 : dirty_0_236; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7243 = 3'h5 == state ? _GEN_6698 : dirty_0_237; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7244 = 3'h5 == state ? _GEN_6699 : dirty_0_238; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7245 = 3'h5 == state ? _GEN_6700 : dirty_0_239; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7246 = 3'h5 == state ? _GEN_6701 : dirty_0_240; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7247 = 3'h5 == state ? _GEN_6702 : dirty_0_241; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7248 = 3'h5 == state ? _GEN_6703 : dirty_0_242; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7249 = 3'h5 == state ? _GEN_6704 : dirty_0_243; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7250 = 3'h5 == state ? _GEN_6705 : dirty_0_244; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7251 = 3'h5 == state ? _GEN_6706 : dirty_0_245; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7252 = 3'h5 == state ? _GEN_6707 : dirty_0_246; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7253 = 3'h5 == state ? _GEN_6708 : dirty_0_247; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7254 = 3'h5 == state ? _GEN_6709 : dirty_0_248; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7255 = 3'h5 == state ? _GEN_6710 : dirty_0_249; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7256 = 3'h5 == state ? _GEN_6711 : dirty_0_250; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7257 = 3'h5 == state ? _GEN_6712 : dirty_0_251; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7258 = 3'h5 == state ? _GEN_6713 : dirty_0_252; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7259 = 3'h5 == state ? _GEN_6714 : dirty_0_253; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7260 = 3'h5 == state ? _GEN_6715 : dirty_0_254; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7261 = 3'h5 == state ? _GEN_6716 : dirty_0_255; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7262 = 3'h5 == state ? _GEN_6717 : dirty_1_0; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7263 = 3'h5 == state ? _GEN_6718 : dirty_1_1; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7264 = 3'h5 == state ? _GEN_6719 : dirty_1_2; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7265 = 3'h5 == state ? _GEN_6720 : dirty_1_3; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7266 = 3'h5 == state ? _GEN_6721 : dirty_1_4; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7267 = 3'h5 == state ? _GEN_6722 : dirty_1_5; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7268 = 3'h5 == state ? _GEN_6723 : dirty_1_6; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7269 = 3'h5 == state ? _GEN_6724 : dirty_1_7; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7270 = 3'h5 == state ? _GEN_6725 : dirty_1_8; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7271 = 3'h5 == state ? _GEN_6726 : dirty_1_9; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7272 = 3'h5 == state ? _GEN_6727 : dirty_1_10; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7273 = 3'h5 == state ? _GEN_6728 : dirty_1_11; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7274 = 3'h5 == state ? _GEN_6729 : dirty_1_12; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7275 = 3'h5 == state ? _GEN_6730 : dirty_1_13; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7276 = 3'h5 == state ? _GEN_6731 : dirty_1_14; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7277 = 3'h5 == state ? _GEN_6732 : dirty_1_15; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7278 = 3'h5 == state ? _GEN_6733 : dirty_1_16; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7279 = 3'h5 == state ? _GEN_6734 : dirty_1_17; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7280 = 3'h5 == state ? _GEN_6735 : dirty_1_18; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7281 = 3'h5 == state ? _GEN_6736 : dirty_1_19; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7282 = 3'h5 == state ? _GEN_6737 : dirty_1_20; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7283 = 3'h5 == state ? _GEN_6738 : dirty_1_21; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7284 = 3'h5 == state ? _GEN_6739 : dirty_1_22; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7285 = 3'h5 == state ? _GEN_6740 : dirty_1_23; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7286 = 3'h5 == state ? _GEN_6741 : dirty_1_24; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7287 = 3'h5 == state ? _GEN_6742 : dirty_1_25; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7288 = 3'h5 == state ? _GEN_6743 : dirty_1_26; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7289 = 3'h5 == state ? _GEN_6744 : dirty_1_27; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7290 = 3'h5 == state ? _GEN_6745 : dirty_1_28; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7291 = 3'h5 == state ? _GEN_6746 : dirty_1_29; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7292 = 3'h5 == state ? _GEN_6747 : dirty_1_30; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7293 = 3'h5 == state ? _GEN_6748 : dirty_1_31; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7294 = 3'h5 == state ? _GEN_6749 : dirty_1_32; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7295 = 3'h5 == state ? _GEN_6750 : dirty_1_33; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7296 = 3'h5 == state ? _GEN_6751 : dirty_1_34; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7297 = 3'h5 == state ? _GEN_6752 : dirty_1_35; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7298 = 3'h5 == state ? _GEN_6753 : dirty_1_36; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7299 = 3'h5 == state ? _GEN_6754 : dirty_1_37; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7300 = 3'h5 == state ? _GEN_6755 : dirty_1_38; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7301 = 3'h5 == state ? _GEN_6756 : dirty_1_39; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7302 = 3'h5 == state ? _GEN_6757 : dirty_1_40; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7303 = 3'h5 == state ? _GEN_6758 : dirty_1_41; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7304 = 3'h5 == state ? _GEN_6759 : dirty_1_42; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7305 = 3'h5 == state ? _GEN_6760 : dirty_1_43; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7306 = 3'h5 == state ? _GEN_6761 : dirty_1_44; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7307 = 3'h5 == state ? _GEN_6762 : dirty_1_45; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7308 = 3'h5 == state ? _GEN_6763 : dirty_1_46; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7309 = 3'h5 == state ? _GEN_6764 : dirty_1_47; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7310 = 3'h5 == state ? _GEN_6765 : dirty_1_48; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7311 = 3'h5 == state ? _GEN_6766 : dirty_1_49; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7312 = 3'h5 == state ? _GEN_6767 : dirty_1_50; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7313 = 3'h5 == state ? _GEN_6768 : dirty_1_51; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7314 = 3'h5 == state ? _GEN_6769 : dirty_1_52; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7315 = 3'h5 == state ? _GEN_6770 : dirty_1_53; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7316 = 3'h5 == state ? _GEN_6771 : dirty_1_54; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7317 = 3'h5 == state ? _GEN_6772 : dirty_1_55; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7318 = 3'h5 == state ? _GEN_6773 : dirty_1_56; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7319 = 3'h5 == state ? _GEN_6774 : dirty_1_57; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7320 = 3'h5 == state ? _GEN_6775 : dirty_1_58; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7321 = 3'h5 == state ? _GEN_6776 : dirty_1_59; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7322 = 3'h5 == state ? _GEN_6777 : dirty_1_60; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7323 = 3'h5 == state ? _GEN_6778 : dirty_1_61; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7324 = 3'h5 == state ? _GEN_6779 : dirty_1_62; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7325 = 3'h5 == state ? _GEN_6780 : dirty_1_63; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7326 = 3'h5 == state ? _GEN_6781 : dirty_1_64; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7327 = 3'h5 == state ? _GEN_6782 : dirty_1_65; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7328 = 3'h5 == state ? _GEN_6783 : dirty_1_66; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7329 = 3'h5 == state ? _GEN_6784 : dirty_1_67; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7330 = 3'h5 == state ? _GEN_6785 : dirty_1_68; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7331 = 3'h5 == state ? _GEN_6786 : dirty_1_69; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7332 = 3'h5 == state ? _GEN_6787 : dirty_1_70; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7333 = 3'h5 == state ? _GEN_6788 : dirty_1_71; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7334 = 3'h5 == state ? _GEN_6789 : dirty_1_72; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7335 = 3'h5 == state ? _GEN_6790 : dirty_1_73; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7336 = 3'h5 == state ? _GEN_6791 : dirty_1_74; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7337 = 3'h5 == state ? _GEN_6792 : dirty_1_75; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7338 = 3'h5 == state ? _GEN_6793 : dirty_1_76; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7339 = 3'h5 == state ? _GEN_6794 : dirty_1_77; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7340 = 3'h5 == state ? _GEN_6795 : dirty_1_78; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7341 = 3'h5 == state ? _GEN_6796 : dirty_1_79; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7342 = 3'h5 == state ? _GEN_6797 : dirty_1_80; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7343 = 3'h5 == state ? _GEN_6798 : dirty_1_81; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7344 = 3'h5 == state ? _GEN_6799 : dirty_1_82; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7345 = 3'h5 == state ? _GEN_6800 : dirty_1_83; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7346 = 3'h5 == state ? _GEN_6801 : dirty_1_84; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7347 = 3'h5 == state ? _GEN_6802 : dirty_1_85; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7348 = 3'h5 == state ? _GEN_6803 : dirty_1_86; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7349 = 3'h5 == state ? _GEN_6804 : dirty_1_87; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7350 = 3'h5 == state ? _GEN_6805 : dirty_1_88; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7351 = 3'h5 == state ? _GEN_6806 : dirty_1_89; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7352 = 3'h5 == state ? _GEN_6807 : dirty_1_90; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7353 = 3'h5 == state ? _GEN_6808 : dirty_1_91; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7354 = 3'h5 == state ? _GEN_6809 : dirty_1_92; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7355 = 3'h5 == state ? _GEN_6810 : dirty_1_93; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7356 = 3'h5 == state ? _GEN_6811 : dirty_1_94; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7357 = 3'h5 == state ? _GEN_6812 : dirty_1_95; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7358 = 3'h5 == state ? _GEN_6813 : dirty_1_96; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7359 = 3'h5 == state ? _GEN_6814 : dirty_1_97; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7360 = 3'h5 == state ? _GEN_6815 : dirty_1_98; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7361 = 3'h5 == state ? _GEN_6816 : dirty_1_99; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7362 = 3'h5 == state ? _GEN_6817 : dirty_1_100; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7363 = 3'h5 == state ? _GEN_6818 : dirty_1_101; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7364 = 3'h5 == state ? _GEN_6819 : dirty_1_102; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7365 = 3'h5 == state ? _GEN_6820 : dirty_1_103; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7366 = 3'h5 == state ? _GEN_6821 : dirty_1_104; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7367 = 3'h5 == state ? _GEN_6822 : dirty_1_105; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7368 = 3'h5 == state ? _GEN_6823 : dirty_1_106; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7369 = 3'h5 == state ? _GEN_6824 : dirty_1_107; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7370 = 3'h5 == state ? _GEN_6825 : dirty_1_108; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7371 = 3'h5 == state ? _GEN_6826 : dirty_1_109; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7372 = 3'h5 == state ? _GEN_6827 : dirty_1_110; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7373 = 3'h5 == state ? _GEN_6828 : dirty_1_111; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7374 = 3'h5 == state ? _GEN_6829 : dirty_1_112; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7375 = 3'h5 == state ? _GEN_6830 : dirty_1_113; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7376 = 3'h5 == state ? _GEN_6831 : dirty_1_114; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7377 = 3'h5 == state ? _GEN_6832 : dirty_1_115; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7378 = 3'h5 == state ? _GEN_6833 : dirty_1_116; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7379 = 3'h5 == state ? _GEN_6834 : dirty_1_117; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7380 = 3'h5 == state ? _GEN_6835 : dirty_1_118; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7381 = 3'h5 == state ? _GEN_6836 : dirty_1_119; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7382 = 3'h5 == state ? _GEN_6837 : dirty_1_120; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7383 = 3'h5 == state ? _GEN_6838 : dirty_1_121; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7384 = 3'h5 == state ? _GEN_6839 : dirty_1_122; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7385 = 3'h5 == state ? _GEN_6840 : dirty_1_123; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7386 = 3'h5 == state ? _GEN_6841 : dirty_1_124; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7387 = 3'h5 == state ? _GEN_6842 : dirty_1_125; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7388 = 3'h5 == state ? _GEN_6843 : dirty_1_126; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7389 = 3'h5 == state ? _GEN_6844 : dirty_1_127; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7390 = 3'h5 == state ? _GEN_6845 : dirty_1_128; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7391 = 3'h5 == state ? _GEN_6846 : dirty_1_129; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7392 = 3'h5 == state ? _GEN_6847 : dirty_1_130; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7393 = 3'h5 == state ? _GEN_6848 : dirty_1_131; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7394 = 3'h5 == state ? _GEN_6849 : dirty_1_132; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7395 = 3'h5 == state ? _GEN_6850 : dirty_1_133; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7396 = 3'h5 == state ? _GEN_6851 : dirty_1_134; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7397 = 3'h5 == state ? _GEN_6852 : dirty_1_135; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7398 = 3'h5 == state ? _GEN_6853 : dirty_1_136; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7399 = 3'h5 == state ? _GEN_6854 : dirty_1_137; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7400 = 3'h5 == state ? _GEN_6855 : dirty_1_138; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7401 = 3'h5 == state ? _GEN_6856 : dirty_1_139; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7402 = 3'h5 == state ? _GEN_6857 : dirty_1_140; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7403 = 3'h5 == state ? _GEN_6858 : dirty_1_141; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7404 = 3'h5 == state ? _GEN_6859 : dirty_1_142; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7405 = 3'h5 == state ? _GEN_6860 : dirty_1_143; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7406 = 3'h5 == state ? _GEN_6861 : dirty_1_144; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7407 = 3'h5 == state ? _GEN_6862 : dirty_1_145; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7408 = 3'h5 == state ? _GEN_6863 : dirty_1_146; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7409 = 3'h5 == state ? _GEN_6864 : dirty_1_147; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7410 = 3'h5 == state ? _GEN_6865 : dirty_1_148; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7411 = 3'h5 == state ? _GEN_6866 : dirty_1_149; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7412 = 3'h5 == state ? _GEN_6867 : dirty_1_150; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7413 = 3'h5 == state ? _GEN_6868 : dirty_1_151; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7414 = 3'h5 == state ? _GEN_6869 : dirty_1_152; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7415 = 3'h5 == state ? _GEN_6870 : dirty_1_153; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7416 = 3'h5 == state ? _GEN_6871 : dirty_1_154; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7417 = 3'h5 == state ? _GEN_6872 : dirty_1_155; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7418 = 3'h5 == state ? _GEN_6873 : dirty_1_156; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7419 = 3'h5 == state ? _GEN_6874 : dirty_1_157; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7420 = 3'h5 == state ? _GEN_6875 : dirty_1_158; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7421 = 3'h5 == state ? _GEN_6876 : dirty_1_159; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7422 = 3'h5 == state ? _GEN_6877 : dirty_1_160; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7423 = 3'h5 == state ? _GEN_6878 : dirty_1_161; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7424 = 3'h5 == state ? _GEN_6879 : dirty_1_162; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7425 = 3'h5 == state ? _GEN_6880 : dirty_1_163; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7426 = 3'h5 == state ? _GEN_6881 : dirty_1_164; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7427 = 3'h5 == state ? _GEN_6882 : dirty_1_165; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7428 = 3'h5 == state ? _GEN_6883 : dirty_1_166; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7429 = 3'h5 == state ? _GEN_6884 : dirty_1_167; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7430 = 3'h5 == state ? _GEN_6885 : dirty_1_168; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7431 = 3'h5 == state ? _GEN_6886 : dirty_1_169; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7432 = 3'h5 == state ? _GEN_6887 : dirty_1_170; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7433 = 3'h5 == state ? _GEN_6888 : dirty_1_171; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7434 = 3'h5 == state ? _GEN_6889 : dirty_1_172; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7435 = 3'h5 == state ? _GEN_6890 : dirty_1_173; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7436 = 3'h5 == state ? _GEN_6891 : dirty_1_174; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7437 = 3'h5 == state ? _GEN_6892 : dirty_1_175; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7438 = 3'h5 == state ? _GEN_6893 : dirty_1_176; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7439 = 3'h5 == state ? _GEN_6894 : dirty_1_177; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7440 = 3'h5 == state ? _GEN_6895 : dirty_1_178; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7441 = 3'h5 == state ? _GEN_6896 : dirty_1_179; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7442 = 3'h5 == state ? _GEN_6897 : dirty_1_180; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7443 = 3'h5 == state ? _GEN_6898 : dirty_1_181; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7444 = 3'h5 == state ? _GEN_6899 : dirty_1_182; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7445 = 3'h5 == state ? _GEN_6900 : dirty_1_183; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7446 = 3'h5 == state ? _GEN_6901 : dirty_1_184; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7447 = 3'h5 == state ? _GEN_6902 : dirty_1_185; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7448 = 3'h5 == state ? _GEN_6903 : dirty_1_186; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7449 = 3'h5 == state ? _GEN_6904 : dirty_1_187; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7450 = 3'h5 == state ? _GEN_6905 : dirty_1_188; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7451 = 3'h5 == state ? _GEN_6906 : dirty_1_189; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7452 = 3'h5 == state ? _GEN_6907 : dirty_1_190; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7453 = 3'h5 == state ? _GEN_6908 : dirty_1_191; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7454 = 3'h5 == state ? _GEN_6909 : dirty_1_192; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7455 = 3'h5 == state ? _GEN_6910 : dirty_1_193; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7456 = 3'h5 == state ? _GEN_6911 : dirty_1_194; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7457 = 3'h5 == state ? _GEN_6912 : dirty_1_195; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7458 = 3'h5 == state ? _GEN_6913 : dirty_1_196; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7459 = 3'h5 == state ? _GEN_6914 : dirty_1_197; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7460 = 3'h5 == state ? _GEN_6915 : dirty_1_198; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7461 = 3'h5 == state ? _GEN_6916 : dirty_1_199; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7462 = 3'h5 == state ? _GEN_6917 : dirty_1_200; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7463 = 3'h5 == state ? _GEN_6918 : dirty_1_201; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7464 = 3'h5 == state ? _GEN_6919 : dirty_1_202; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7465 = 3'h5 == state ? _GEN_6920 : dirty_1_203; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7466 = 3'h5 == state ? _GEN_6921 : dirty_1_204; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7467 = 3'h5 == state ? _GEN_6922 : dirty_1_205; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7468 = 3'h5 == state ? _GEN_6923 : dirty_1_206; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7469 = 3'h5 == state ? _GEN_6924 : dirty_1_207; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7470 = 3'h5 == state ? _GEN_6925 : dirty_1_208; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7471 = 3'h5 == state ? _GEN_6926 : dirty_1_209; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7472 = 3'h5 == state ? _GEN_6927 : dirty_1_210; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7473 = 3'h5 == state ? _GEN_6928 : dirty_1_211; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7474 = 3'h5 == state ? _GEN_6929 : dirty_1_212; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7475 = 3'h5 == state ? _GEN_6930 : dirty_1_213; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7476 = 3'h5 == state ? _GEN_6931 : dirty_1_214; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7477 = 3'h5 == state ? _GEN_6932 : dirty_1_215; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7478 = 3'h5 == state ? _GEN_6933 : dirty_1_216; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7479 = 3'h5 == state ? _GEN_6934 : dirty_1_217; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7480 = 3'h5 == state ? _GEN_6935 : dirty_1_218; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7481 = 3'h5 == state ? _GEN_6936 : dirty_1_219; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7482 = 3'h5 == state ? _GEN_6937 : dirty_1_220; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7483 = 3'h5 == state ? _GEN_6938 : dirty_1_221; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7484 = 3'h5 == state ? _GEN_6939 : dirty_1_222; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7485 = 3'h5 == state ? _GEN_6940 : dirty_1_223; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7486 = 3'h5 == state ? _GEN_6941 : dirty_1_224; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7487 = 3'h5 == state ? _GEN_6942 : dirty_1_225; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7488 = 3'h5 == state ? _GEN_6943 : dirty_1_226; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7489 = 3'h5 == state ? _GEN_6944 : dirty_1_227; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7490 = 3'h5 == state ? _GEN_6945 : dirty_1_228; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7491 = 3'h5 == state ? _GEN_6946 : dirty_1_229; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7492 = 3'h5 == state ? _GEN_6947 : dirty_1_230; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7493 = 3'h5 == state ? _GEN_6948 : dirty_1_231; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7494 = 3'h5 == state ? _GEN_6949 : dirty_1_232; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7495 = 3'h5 == state ? _GEN_6950 : dirty_1_233; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7496 = 3'h5 == state ? _GEN_6951 : dirty_1_234; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7497 = 3'h5 == state ? _GEN_6952 : dirty_1_235; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7498 = 3'h5 == state ? _GEN_6953 : dirty_1_236; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7499 = 3'h5 == state ? _GEN_6954 : dirty_1_237; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7500 = 3'h5 == state ? _GEN_6955 : dirty_1_238; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7501 = 3'h5 == state ? _GEN_6956 : dirty_1_239; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7502 = 3'h5 == state ? _GEN_6957 : dirty_1_240; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7503 = 3'h5 == state ? _GEN_6958 : dirty_1_241; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7504 = 3'h5 == state ? _GEN_6959 : dirty_1_242; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7505 = 3'h5 == state ? _GEN_6960 : dirty_1_243; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7506 = 3'h5 == state ? _GEN_6961 : dirty_1_244; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7507 = 3'h5 == state ? _GEN_6962 : dirty_1_245; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7508 = 3'h5 == state ? _GEN_6963 : dirty_1_246; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7509 = 3'h5 == state ? _GEN_6964 : dirty_1_247; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7510 = 3'h5 == state ? _GEN_6965 : dirty_1_248; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7511 = 3'h5 == state ? _GEN_6966 : dirty_1_249; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7512 = 3'h5 == state ? _GEN_6967 : dirty_1_250; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7513 = 3'h5 == state ? _GEN_6968 : dirty_1_251; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7514 = 3'h5 == state ? _GEN_6969 : dirty_1_252; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7515 = 3'h5 == state ? _GEN_6970 : dirty_1_253; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7516 = 3'h5 == state ? _GEN_6971 : dirty_1_254; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7517 = 3'h5 == state ? _GEN_6972 : dirty_1_255; // @[dcache.scala 183:18 113:28]
  wire [20:0] _GEN_7520 = 3'h5 == state ? _GEN_6975 : 21'h0; // @[dcache.scala 183:18 143:25]
  wire [20:0] _GEN_7521 = 3'h5 == state ? _GEN_6976 : 21'h0; // @[dcache.scala 183:18 143:25]
  wire [31:0] _GEN_7523 = 3'h5 == state ? _GEN_6978 : 32'h7777; // @[dcache.scala 183:18 155:25]
  wire  _GEN_7524 = 3'h5 == state ? _GEN_6979 : req_valid; // @[dcache.scala 183:18 116:34]
  wire [21:0] _GEN_7526 = 3'h5 == state ? _GEN_6981 : 22'h0; // @[dcache.scala 183:18 98:21]
  wire  _GEN_7527 = 3'h5 == state ? _GEN_6982 : cacheInst_r; // @[dcache.scala 183:18 89:38]
  wire  _GEN_7528 = 3'h5 == state ? _GEN_6983 : invalidate; // @[dcache.scala 183:18 90:38]
  wire  _GEN_7529 = 3'h5 == state ? _GEN_6984 : indexOnly; // @[dcache.scala 183:18 94:38]
  wire  _GEN_7530 = 3'h5 == state ? _GEN_6985 : writeBack; // @[dcache.scala 183:18 93:38]
  wire  _GEN_7531 = 3'h5 == state ? _GEN_6986 : storeTag; // @[dcache.scala 183:18 92:38]
  wire  _GEN_7532 = 3'h5 == state ? _GEN_6987 : loadTag; // @[dcache.scala 183:18 91:38]
  wire [2:0] _GEN_7533 = 3'h4 == state ? _GEN_713 : _GEN_6988; // @[dcache.scala 183:18]
  wire [2:0] _GEN_7535 = 3'h4 == state ? _GEN_715 : 3'h0; // @[dcache.scala 183:18 159:25]
  wire [31:0] _GEN_7536 = 3'h4 == state ? _GEN_716 : 32'h0; // @[dcache.scala 183:18 160:25]
  wire [1:0] _GEN_7537 = 3'h4 == state ? wr_cnt : _GEN_6989; // @[dcache.scala 183:18 178:34]
  wire [31:0] _GEN_7538 = 3'h4 == state ? 32'h0 : _GEN_6990; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_7539 = 3'h4 == state ? 32'h0 : _GEN_6991; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_7540 = 3'h4 == state ? 32'h0 : _GEN_6992; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_7541 = 3'h4 == state ? 32'h0 : _GEN_6993; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_7542 = 3'h4 == state ? 32'h0 : _GEN_6994; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_7543 = 3'h4 == state ? 32'h0 : _GEN_6995; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_7544 = 3'h4 == state ? 32'h0 : _GEN_6996; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_7545 = 3'h4 == state ? 32'h0 : _GEN_6997; // @[dcache.scala 183:18 149:33]
  wire [3:0] _GEN_7546 = 3'h4 == state ? 4'h0 : _GEN_6998; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7547 = 3'h4 == state ? 4'h0 : _GEN_6999; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7548 = 3'h4 == state ? 4'h0 : _GEN_7000; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7549 = 3'h4 == state ? 4'h0 : _GEN_7001; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7550 = 3'h4 == state ? 4'h0 : _GEN_7002; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7551 = 3'h4 == state ? 4'h0 : _GEN_7003; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7552 = 3'h4 == state ? 4'h0 : _GEN_7004; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_7553 = 3'h4 == state ? 4'h0 : _GEN_7005; // @[dcache.scala 183:18 150:33]
  wire  _GEN_7554 = 3'h4 == state ? dirty_0_0 : _GEN_7006; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7555 = 3'h4 == state ? dirty_0_1 : _GEN_7007; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7556 = 3'h4 == state ? dirty_0_2 : _GEN_7008; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7557 = 3'h4 == state ? dirty_0_3 : _GEN_7009; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7558 = 3'h4 == state ? dirty_0_4 : _GEN_7010; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7559 = 3'h4 == state ? dirty_0_5 : _GEN_7011; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7560 = 3'h4 == state ? dirty_0_6 : _GEN_7012; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7561 = 3'h4 == state ? dirty_0_7 : _GEN_7013; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7562 = 3'h4 == state ? dirty_0_8 : _GEN_7014; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7563 = 3'h4 == state ? dirty_0_9 : _GEN_7015; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7564 = 3'h4 == state ? dirty_0_10 : _GEN_7016; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7565 = 3'h4 == state ? dirty_0_11 : _GEN_7017; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7566 = 3'h4 == state ? dirty_0_12 : _GEN_7018; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7567 = 3'h4 == state ? dirty_0_13 : _GEN_7019; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7568 = 3'h4 == state ? dirty_0_14 : _GEN_7020; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7569 = 3'h4 == state ? dirty_0_15 : _GEN_7021; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7570 = 3'h4 == state ? dirty_0_16 : _GEN_7022; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7571 = 3'h4 == state ? dirty_0_17 : _GEN_7023; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7572 = 3'h4 == state ? dirty_0_18 : _GEN_7024; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7573 = 3'h4 == state ? dirty_0_19 : _GEN_7025; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7574 = 3'h4 == state ? dirty_0_20 : _GEN_7026; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7575 = 3'h4 == state ? dirty_0_21 : _GEN_7027; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7576 = 3'h4 == state ? dirty_0_22 : _GEN_7028; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7577 = 3'h4 == state ? dirty_0_23 : _GEN_7029; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7578 = 3'h4 == state ? dirty_0_24 : _GEN_7030; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7579 = 3'h4 == state ? dirty_0_25 : _GEN_7031; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7580 = 3'h4 == state ? dirty_0_26 : _GEN_7032; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7581 = 3'h4 == state ? dirty_0_27 : _GEN_7033; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7582 = 3'h4 == state ? dirty_0_28 : _GEN_7034; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7583 = 3'h4 == state ? dirty_0_29 : _GEN_7035; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7584 = 3'h4 == state ? dirty_0_30 : _GEN_7036; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7585 = 3'h4 == state ? dirty_0_31 : _GEN_7037; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7586 = 3'h4 == state ? dirty_0_32 : _GEN_7038; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7587 = 3'h4 == state ? dirty_0_33 : _GEN_7039; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7588 = 3'h4 == state ? dirty_0_34 : _GEN_7040; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7589 = 3'h4 == state ? dirty_0_35 : _GEN_7041; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7590 = 3'h4 == state ? dirty_0_36 : _GEN_7042; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7591 = 3'h4 == state ? dirty_0_37 : _GEN_7043; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7592 = 3'h4 == state ? dirty_0_38 : _GEN_7044; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7593 = 3'h4 == state ? dirty_0_39 : _GEN_7045; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7594 = 3'h4 == state ? dirty_0_40 : _GEN_7046; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7595 = 3'h4 == state ? dirty_0_41 : _GEN_7047; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7596 = 3'h4 == state ? dirty_0_42 : _GEN_7048; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7597 = 3'h4 == state ? dirty_0_43 : _GEN_7049; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7598 = 3'h4 == state ? dirty_0_44 : _GEN_7050; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7599 = 3'h4 == state ? dirty_0_45 : _GEN_7051; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7600 = 3'h4 == state ? dirty_0_46 : _GEN_7052; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7601 = 3'h4 == state ? dirty_0_47 : _GEN_7053; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7602 = 3'h4 == state ? dirty_0_48 : _GEN_7054; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7603 = 3'h4 == state ? dirty_0_49 : _GEN_7055; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7604 = 3'h4 == state ? dirty_0_50 : _GEN_7056; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7605 = 3'h4 == state ? dirty_0_51 : _GEN_7057; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7606 = 3'h4 == state ? dirty_0_52 : _GEN_7058; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7607 = 3'h4 == state ? dirty_0_53 : _GEN_7059; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7608 = 3'h4 == state ? dirty_0_54 : _GEN_7060; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7609 = 3'h4 == state ? dirty_0_55 : _GEN_7061; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7610 = 3'h4 == state ? dirty_0_56 : _GEN_7062; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7611 = 3'h4 == state ? dirty_0_57 : _GEN_7063; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7612 = 3'h4 == state ? dirty_0_58 : _GEN_7064; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7613 = 3'h4 == state ? dirty_0_59 : _GEN_7065; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7614 = 3'h4 == state ? dirty_0_60 : _GEN_7066; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7615 = 3'h4 == state ? dirty_0_61 : _GEN_7067; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7616 = 3'h4 == state ? dirty_0_62 : _GEN_7068; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7617 = 3'h4 == state ? dirty_0_63 : _GEN_7069; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7618 = 3'h4 == state ? dirty_0_64 : _GEN_7070; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7619 = 3'h4 == state ? dirty_0_65 : _GEN_7071; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7620 = 3'h4 == state ? dirty_0_66 : _GEN_7072; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7621 = 3'h4 == state ? dirty_0_67 : _GEN_7073; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7622 = 3'h4 == state ? dirty_0_68 : _GEN_7074; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7623 = 3'h4 == state ? dirty_0_69 : _GEN_7075; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7624 = 3'h4 == state ? dirty_0_70 : _GEN_7076; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7625 = 3'h4 == state ? dirty_0_71 : _GEN_7077; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7626 = 3'h4 == state ? dirty_0_72 : _GEN_7078; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7627 = 3'h4 == state ? dirty_0_73 : _GEN_7079; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7628 = 3'h4 == state ? dirty_0_74 : _GEN_7080; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7629 = 3'h4 == state ? dirty_0_75 : _GEN_7081; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7630 = 3'h4 == state ? dirty_0_76 : _GEN_7082; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7631 = 3'h4 == state ? dirty_0_77 : _GEN_7083; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7632 = 3'h4 == state ? dirty_0_78 : _GEN_7084; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7633 = 3'h4 == state ? dirty_0_79 : _GEN_7085; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7634 = 3'h4 == state ? dirty_0_80 : _GEN_7086; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7635 = 3'h4 == state ? dirty_0_81 : _GEN_7087; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7636 = 3'h4 == state ? dirty_0_82 : _GEN_7088; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7637 = 3'h4 == state ? dirty_0_83 : _GEN_7089; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7638 = 3'h4 == state ? dirty_0_84 : _GEN_7090; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7639 = 3'h4 == state ? dirty_0_85 : _GEN_7091; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7640 = 3'h4 == state ? dirty_0_86 : _GEN_7092; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7641 = 3'h4 == state ? dirty_0_87 : _GEN_7093; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7642 = 3'h4 == state ? dirty_0_88 : _GEN_7094; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7643 = 3'h4 == state ? dirty_0_89 : _GEN_7095; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7644 = 3'h4 == state ? dirty_0_90 : _GEN_7096; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7645 = 3'h4 == state ? dirty_0_91 : _GEN_7097; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7646 = 3'h4 == state ? dirty_0_92 : _GEN_7098; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7647 = 3'h4 == state ? dirty_0_93 : _GEN_7099; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7648 = 3'h4 == state ? dirty_0_94 : _GEN_7100; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7649 = 3'h4 == state ? dirty_0_95 : _GEN_7101; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7650 = 3'h4 == state ? dirty_0_96 : _GEN_7102; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7651 = 3'h4 == state ? dirty_0_97 : _GEN_7103; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7652 = 3'h4 == state ? dirty_0_98 : _GEN_7104; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7653 = 3'h4 == state ? dirty_0_99 : _GEN_7105; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7654 = 3'h4 == state ? dirty_0_100 : _GEN_7106; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7655 = 3'h4 == state ? dirty_0_101 : _GEN_7107; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7656 = 3'h4 == state ? dirty_0_102 : _GEN_7108; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7657 = 3'h4 == state ? dirty_0_103 : _GEN_7109; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7658 = 3'h4 == state ? dirty_0_104 : _GEN_7110; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7659 = 3'h4 == state ? dirty_0_105 : _GEN_7111; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7660 = 3'h4 == state ? dirty_0_106 : _GEN_7112; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7661 = 3'h4 == state ? dirty_0_107 : _GEN_7113; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7662 = 3'h4 == state ? dirty_0_108 : _GEN_7114; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7663 = 3'h4 == state ? dirty_0_109 : _GEN_7115; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7664 = 3'h4 == state ? dirty_0_110 : _GEN_7116; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7665 = 3'h4 == state ? dirty_0_111 : _GEN_7117; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7666 = 3'h4 == state ? dirty_0_112 : _GEN_7118; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7667 = 3'h4 == state ? dirty_0_113 : _GEN_7119; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7668 = 3'h4 == state ? dirty_0_114 : _GEN_7120; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7669 = 3'h4 == state ? dirty_0_115 : _GEN_7121; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7670 = 3'h4 == state ? dirty_0_116 : _GEN_7122; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7671 = 3'h4 == state ? dirty_0_117 : _GEN_7123; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7672 = 3'h4 == state ? dirty_0_118 : _GEN_7124; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7673 = 3'h4 == state ? dirty_0_119 : _GEN_7125; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7674 = 3'h4 == state ? dirty_0_120 : _GEN_7126; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7675 = 3'h4 == state ? dirty_0_121 : _GEN_7127; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7676 = 3'h4 == state ? dirty_0_122 : _GEN_7128; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7677 = 3'h4 == state ? dirty_0_123 : _GEN_7129; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7678 = 3'h4 == state ? dirty_0_124 : _GEN_7130; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7679 = 3'h4 == state ? dirty_0_125 : _GEN_7131; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7680 = 3'h4 == state ? dirty_0_126 : _GEN_7132; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7681 = 3'h4 == state ? dirty_0_127 : _GEN_7133; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7682 = 3'h4 == state ? dirty_0_128 : _GEN_7134; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7683 = 3'h4 == state ? dirty_0_129 : _GEN_7135; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7684 = 3'h4 == state ? dirty_0_130 : _GEN_7136; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7685 = 3'h4 == state ? dirty_0_131 : _GEN_7137; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7686 = 3'h4 == state ? dirty_0_132 : _GEN_7138; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7687 = 3'h4 == state ? dirty_0_133 : _GEN_7139; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7688 = 3'h4 == state ? dirty_0_134 : _GEN_7140; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7689 = 3'h4 == state ? dirty_0_135 : _GEN_7141; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7690 = 3'h4 == state ? dirty_0_136 : _GEN_7142; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7691 = 3'h4 == state ? dirty_0_137 : _GEN_7143; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7692 = 3'h4 == state ? dirty_0_138 : _GEN_7144; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7693 = 3'h4 == state ? dirty_0_139 : _GEN_7145; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7694 = 3'h4 == state ? dirty_0_140 : _GEN_7146; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7695 = 3'h4 == state ? dirty_0_141 : _GEN_7147; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7696 = 3'h4 == state ? dirty_0_142 : _GEN_7148; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7697 = 3'h4 == state ? dirty_0_143 : _GEN_7149; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7698 = 3'h4 == state ? dirty_0_144 : _GEN_7150; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7699 = 3'h4 == state ? dirty_0_145 : _GEN_7151; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7700 = 3'h4 == state ? dirty_0_146 : _GEN_7152; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7701 = 3'h4 == state ? dirty_0_147 : _GEN_7153; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7702 = 3'h4 == state ? dirty_0_148 : _GEN_7154; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7703 = 3'h4 == state ? dirty_0_149 : _GEN_7155; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7704 = 3'h4 == state ? dirty_0_150 : _GEN_7156; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7705 = 3'h4 == state ? dirty_0_151 : _GEN_7157; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7706 = 3'h4 == state ? dirty_0_152 : _GEN_7158; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7707 = 3'h4 == state ? dirty_0_153 : _GEN_7159; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7708 = 3'h4 == state ? dirty_0_154 : _GEN_7160; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7709 = 3'h4 == state ? dirty_0_155 : _GEN_7161; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7710 = 3'h4 == state ? dirty_0_156 : _GEN_7162; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7711 = 3'h4 == state ? dirty_0_157 : _GEN_7163; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7712 = 3'h4 == state ? dirty_0_158 : _GEN_7164; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7713 = 3'h4 == state ? dirty_0_159 : _GEN_7165; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7714 = 3'h4 == state ? dirty_0_160 : _GEN_7166; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7715 = 3'h4 == state ? dirty_0_161 : _GEN_7167; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7716 = 3'h4 == state ? dirty_0_162 : _GEN_7168; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7717 = 3'h4 == state ? dirty_0_163 : _GEN_7169; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7718 = 3'h4 == state ? dirty_0_164 : _GEN_7170; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7719 = 3'h4 == state ? dirty_0_165 : _GEN_7171; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7720 = 3'h4 == state ? dirty_0_166 : _GEN_7172; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7721 = 3'h4 == state ? dirty_0_167 : _GEN_7173; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7722 = 3'h4 == state ? dirty_0_168 : _GEN_7174; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7723 = 3'h4 == state ? dirty_0_169 : _GEN_7175; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7724 = 3'h4 == state ? dirty_0_170 : _GEN_7176; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7725 = 3'h4 == state ? dirty_0_171 : _GEN_7177; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7726 = 3'h4 == state ? dirty_0_172 : _GEN_7178; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7727 = 3'h4 == state ? dirty_0_173 : _GEN_7179; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7728 = 3'h4 == state ? dirty_0_174 : _GEN_7180; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7729 = 3'h4 == state ? dirty_0_175 : _GEN_7181; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7730 = 3'h4 == state ? dirty_0_176 : _GEN_7182; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7731 = 3'h4 == state ? dirty_0_177 : _GEN_7183; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7732 = 3'h4 == state ? dirty_0_178 : _GEN_7184; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7733 = 3'h4 == state ? dirty_0_179 : _GEN_7185; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7734 = 3'h4 == state ? dirty_0_180 : _GEN_7186; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7735 = 3'h4 == state ? dirty_0_181 : _GEN_7187; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7736 = 3'h4 == state ? dirty_0_182 : _GEN_7188; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7737 = 3'h4 == state ? dirty_0_183 : _GEN_7189; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7738 = 3'h4 == state ? dirty_0_184 : _GEN_7190; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7739 = 3'h4 == state ? dirty_0_185 : _GEN_7191; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7740 = 3'h4 == state ? dirty_0_186 : _GEN_7192; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7741 = 3'h4 == state ? dirty_0_187 : _GEN_7193; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7742 = 3'h4 == state ? dirty_0_188 : _GEN_7194; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7743 = 3'h4 == state ? dirty_0_189 : _GEN_7195; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7744 = 3'h4 == state ? dirty_0_190 : _GEN_7196; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7745 = 3'h4 == state ? dirty_0_191 : _GEN_7197; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7746 = 3'h4 == state ? dirty_0_192 : _GEN_7198; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7747 = 3'h4 == state ? dirty_0_193 : _GEN_7199; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7748 = 3'h4 == state ? dirty_0_194 : _GEN_7200; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7749 = 3'h4 == state ? dirty_0_195 : _GEN_7201; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7750 = 3'h4 == state ? dirty_0_196 : _GEN_7202; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7751 = 3'h4 == state ? dirty_0_197 : _GEN_7203; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7752 = 3'h4 == state ? dirty_0_198 : _GEN_7204; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7753 = 3'h4 == state ? dirty_0_199 : _GEN_7205; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7754 = 3'h4 == state ? dirty_0_200 : _GEN_7206; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7755 = 3'h4 == state ? dirty_0_201 : _GEN_7207; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7756 = 3'h4 == state ? dirty_0_202 : _GEN_7208; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7757 = 3'h4 == state ? dirty_0_203 : _GEN_7209; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7758 = 3'h4 == state ? dirty_0_204 : _GEN_7210; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7759 = 3'h4 == state ? dirty_0_205 : _GEN_7211; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7760 = 3'h4 == state ? dirty_0_206 : _GEN_7212; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7761 = 3'h4 == state ? dirty_0_207 : _GEN_7213; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7762 = 3'h4 == state ? dirty_0_208 : _GEN_7214; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7763 = 3'h4 == state ? dirty_0_209 : _GEN_7215; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7764 = 3'h4 == state ? dirty_0_210 : _GEN_7216; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7765 = 3'h4 == state ? dirty_0_211 : _GEN_7217; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7766 = 3'h4 == state ? dirty_0_212 : _GEN_7218; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7767 = 3'h4 == state ? dirty_0_213 : _GEN_7219; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7768 = 3'h4 == state ? dirty_0_214 : _GEN_7220; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7769 = 3'h4 == state ? dirty_0_215 : _GEN_7221; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7770 = 3'h4 == state ? dirty_0_216 : _GEN_7222; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7771 = 3'h4 == state ? dirty_0_217 : _GEN_7223; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7772 = 3'h4 == state ? dirty_0_218 : _GEN_7224; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7773 = 3'h4 == state ? dirty_0_219 : _GEN_7225; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7774 = 3'h4 == state ? dirty_0_220 : _GEN_7226; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7775 = 3'h4 == state ? dirty_0_221 : _GEN_7227; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7776 = 3'h4 == state ? dirty_0_222 : _GEN_7228; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7777 = 3'h4 == state ? dirty_0_223 : _GEN_7229; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7778 = 3'h4 == state ? dirty_0_224 : _GEN_7230; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7779 = 3'h4 == state ? dirty_0_225 : _GEN_7231; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7780 = 3'h4 == state ? dirty_0_226 : _GEN_7232; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7781 = 3'h4 == state ? dirty_0_227 : _GEN_7233; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7782 = 3'h4 == state ? dirty_0_228 : _GEN_7234; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7783 = 3'h4 == state ? dirty_0_229 : _GEN_7235; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7784 = 3'h4 == state ? dirty_0_230 : _GEN_7236; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7785 = 3'h4 == state ? dirty_0_231 : _GEN_7237; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7786 = 3'h4 == state ? dirty_0_232 : _GEN_7238; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7787 = 3'h4 == state ? dirty_0_233 : _GEN_7239; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7788 = 3'h4 == state ? dirty_0_234 : _GEN_7240; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7789 = 3'h4 == state ? dirty_0_235 : _GEN_7241; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7790 = 3'h4 == state ? dirty_0_236 : _GEN_7242; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7791 = 3'h4 == state ? dirty_0_237 : _GEN_7243; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7792 = 3'h4 == state ? dirty_0_238 : _GEN_7244; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7793 = 3'h4 == state ? dirty_0_239 : _GEN_7245; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7794 = 3'h4 == state ? dirty_0_240 : _GEN_7246; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7795 = 3'h4 == state ? dirty_0_241 : _GEN_7247; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7796 = 3'h4 == state ? dirty_0_242 : _GEN_7248; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7797 = 3'h4 == state ? dirty_0_243 : _GEN_7249; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7798 = 3'h4 == state ? dirty_0_244 : _GEN_7250; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7799 = 3'h4 == state ? dirty_0_245 : _GEN_7251; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7800 = 3'h4 == state ? dirty_0_246 : _GEN_7252; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7801 = 3'h4 == state ? dirty_0_247 : _GEN_7253; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7802 = 3'h4 == state ? dirty_0_248 : _GEN_7254; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7803 = 3'h4 == state ? dirty_0_249 : _GEN_7255; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7804 = 3'h4 == state ? dirty_0_250 : _GEN_7256; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7805 = 3'h4 == state ? dirty_0_251 : _GEN_7257; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7806 = 3'h4 == state ? dirty_0_252 : _GEN_7258; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7807 = 3'h4 == state ? dirty_0_253 : _GEN_7259; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7808 = 3'h4 == state ? dirty_0_254 : _GEN_7260; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7809 = 3'h4 == state ? dirty_0_255 : _GEN_7261; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7810 = 3'h4 == state ? dirty_1_0 : _GEN_7262; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7811 = 3'h4 == state ? dirty_1_1 : _GEN_7263; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7812 = 3'h4 == state ? dirty_1_2 : _GEN_7264; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7813 = 3'h4 == state ? dirty_1_3 : _GEN_7265; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7814 = 3'h4 == state ? dirty_1_4 : _GEN_7266; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7815 = 3'h4 == state ? dirty_1_5 : _GEN_7267; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7816 = 3'h4 == state ? dirty_1_6 : _GEN_7268; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7817 = 3'h4 == state ? dirty_1_7 : _GEN_7269; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7818 = 3'h4 == state ? dirty_1_8 : _GEN_7270; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7819 = 3'h4 == state ? dirty_1_9 : _GEN_7271; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7820 = 3'h4 == state ? dirty_1_10 : _GEN_7272; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7821 = 3'h4 == state ? dirty_1_11 : _GEN_7273; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7822 = 3'h4 == state ? dirty_1_12 : _GEN_7274; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7823 = 3'h4 == state ? dirty_1_13 : _GEN_7275; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7824 = 3'h4 == state ? dirty_1_14 : _GEN_7276; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7825 = 3'h4 == state ? dirty_1_15 : _GEN_7277; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7826 = 3'h4 == state ? dirty_1_16 : _GEN_7278; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7827 = 3'h4 == state ? dirty_1_17 : _GEN_7279; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7828 = 3'h4 == state ? dirty_1_18 : _GEN_7280; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7829 = 3'h4 == state ? dirty_1_19 : _GEN_7281; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7830 = 3'h4 == state ? dirty_1_20 : _GEN_7282; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7831 = 3'h4 == state ? dirty_1_21 : _GEN_7283; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7832 = 3'h4 == state ? dirty_1_22 : _GEN_7284; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7833 = 3'h4 == state ? dirty_1_23 : _GEN_7285; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7834 = 3'h4 == state ? dirty_1_24 : _GEN_7286; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7835 = 3'h4 == state ? dirty_1_25 : _GEN_7287; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7836 = 3'h4 == state ? dirty_1_26 : _GEN_7288; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7837 = 3'h4 == state ? dirty_1_27 : _GEN_7289; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7838 = 3'h4 == state ? dirty_1_28 : _GEN_7290; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7839 = 3'h4 == state ? dirty_1_29 : _GEN_7291; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7840 = 3'h4 == state ? dirty_1_30 : _GEN_7292; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7841 = 3'h4 == state ? dirty_1_31 : _GEN_7293; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7842 = 3'h4 == state ? dirty_1_32 : _GEN_7294; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7843 = 3'h4 == state ? dirty_1_33 : _GEN_7295; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7844 = 3'h4 == state ? dirty_1_34 : _GEN_7296; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7845 = 3'h4 == state ? dirty_1_35 : _GEN_7297; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7846 = 3'h4 == state ? dirty_1_36 : _GEN_7298; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7847 = 3'h4 == state ? dirty_1_37 : _GEN_7299; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7848 = 3'h4 == state ? dirty_1_38 : _GEN_7300; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7849 = 3'h4 == state ? dirty_1_39 : _GEN_7301; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7850 = 3'h4 == state ? dirty_1_40 : _GEN_7302; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7851 = 3'h4 == state ? dirty_1_41 : _GEN_7303; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7852 = 3'h4 == state ? dirty_1_42 : _GEN_7304; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7853 = 3'h4 == state ? dirty_1_43 : _GEN_7305; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7854 = 3'h4 == state ? dirty_1_44 : _GEN_7306; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7855 = 3'h4 == state ? dirty_1_45 : _GEN_7307; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7856 = 3'h4 == state ? dirty_1_46 : _GEN_7308; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7857 = 3'h4 == state ? dirty_1_47 : _GEN_7309; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7858 = 3'h4 == state ? dirty_1_48 : _GEN_7310; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7859 = 3'h4 == state ? dirty_1_49 : _GEN_7311; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7860 = 3'h4 == state ? dirty_1_50 : _GEN_7312; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7861 = 3'h4 == state ? dirty_1_51 : _GEN_7313; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7862 = 3'h4 == state ? dirty_1_52 : _GEN_7314; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7863 = 3'h4 == state ? dirty_1_53 : _GEN_7315; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7864 = 3'h4 == state ? dirty_1_54 : _GEN_7316; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7865 = 3'h4 == state ? dirty_1_55 : _GEN_7317; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7866 = 3'h4 == state ? dirty_1_56 : _GEN_7318; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7867 = 3'h4 == state ? dirty_1_57 : _GEN_7319; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7868 = 3'h4 == state ? dirty_1_58 : _GEN_7320; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7869 = 3'h4 == state ? dirty_1_59 : _GEN_7321; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7870 = 3'h4 == state ? dirty_1_60 : _GEN_7322; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7871 = 3'h4 == state ? dirty_1_61 : _GEN_7323; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7872 = 3'h4 == state ? dirty_1_62 : _GEN_7324; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7873 = 3'h4 == state ? dirty_1_63 : _GEN_7325; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7874 = 3'h4 == state ? dirty_1_64 : _GEN_7326; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7875 = 3'h4 == state ? dirty_1_65 : _GEN_7327; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7876 = 3'h4 == state ? dirty_1_66 : _GEN_7328; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7877 = 3'h4 == state ? dirty_1_67 : _GEN_7329; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7878 = 3'h4 == state ? dirty_1_68 : _GEN_7330; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7879 = 3'h4 == state ? dirty_1_69 : _GEN_7331; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7880 = 3'h4 == state ? dirty_1_70 : _GEN_7332; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7881 = 3'h4 == state ? dirty_1_71 : _GEN_7333; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7882 = 3'h4 == state ? dirty_1_72 : _GEN_7334; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7883 = 3'h4 == state ? dirty_1_73 : _GEN_7335; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7884 = 3'h4 == state ? dirty_1_74 : _GEN_7336; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7885 = 3'h4 == state ? dirty_1_75 : _GEN_7337; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7886 = 3'h4 == state ? dirty_1_76 : _GEN_7338; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7887 = 3'h4 == state ? dirty_1_77 : _GEN_7339; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7888 = 3'h4 == state ? dirty_1_78 : _GEN_7340; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7889 = 3'h4 == state ? dirty_1_79 : _GEN_7341; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7890 = 3'h4 == state ? dirty_1_80 : _GEN_7342; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7891 = 3'h4 == state ? dirty_1_81 : _GEN_7343; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7892 = 3'h4 == state ? dirty_1_82 : _GEN_7344; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7893 = 3'h4 == state ? dirty_1_83 : _GEN_7345; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7894 = 3'h4 == state ? dirty_1_84 : _GEN_7346; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7895 = 3'h4 == state ? dirty_1_85 : _GEN_7347; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7896 = 3'h4 == state ? dirty_1_86 : _GEN_7348; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7897 = 3'h4 == state ? dirty_1_87 : _GEN_7349; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7898 = 3'h4 == state ? dirty_1_88 : _GEN_7350; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7899 = 3'h4 == state ? dirty_1_89 : _GEN_7351; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7900 = 3'h4 == state ? dirty_1_90 : _GEN_7352; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7901 = 3'h4 == state ? dirty_1_91 : _GEN_7353; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7902 = 3'h4 == state ? dirty_1_92 : _GEN_7354; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7903 = 3'h4 == state ? dirty_1_93 : _GEN_7355; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7904 = 3'h4 == state ? dirty_1_94 : _GEN_7356; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7905 = 3'h4 == state ? dirty_1_95 : _GEN_7357; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7906 = 3'h4 == state ? dirty_1_96 : _GEN_7358; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7907 = 3'h4 == state ? dirty_1_97 : _GEN_7359; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7908 = 3'h4 == state ? dirty_1_98 : _GEN_7360; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7909 = 3'h4 == state ? dirty_1_99 : _GEN_7361; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7910 = 3'h4 == state ? dirty_1_100 : _GEN_7362; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7911 = 3'h4 == state ? dirty_1_101 : _GEN_7363; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7912 = 3'h4 == state ? dirty_1_102 : _GEN_7364; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7913 = 3'h4 == state ? dirty_1_103 : _GEN_7365; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7914 = 3'h4 == state ? dirty_1_104 : _GEN_7366; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7915 = 3'h4 == state ? dirty_1_105 : _GEN_7367; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7916 = 3'h4 == state ? dirty_1_106 : _GEN_7368; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7917 = 3'h4 == state ? dirty_1_107 : _GEN_7369; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7918 = 3'h4 == state ? dirty_1_108 : _GEN_7370; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7919 = 3'h4 == state ? dirty_1_109 : _GEN_7371; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7920 = 3'h4 == state ? dirty_1_110 : _GEN_7372; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7921 = 3'h4 == state ? dirty_1_111 : _GEN_7373; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7922 = 3'h4 == state ? dirty_1_112 : _GEN_7374; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7923 = 3'h4 == state ? dirty_1_113 : _GEN_7375; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7924 = 3'h4 == state ? dirty_1_114 : _GEN_7376; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7925 = 3'h4 == state ? dirty_1_115 : _GEN_7377; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7926 = 3'h4 == state ? dirty_1_116 : _GEN_7378; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7927 = 3'h4 == state ? dirty_1_117 : _GEN_7379; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7928 = 3'h4 == state ? dirty_1_118 : _GEN_7380; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7929 = 3'h4 == state ? dirty_1_119 : _GEN_7381; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7930 = 3'h4 == state ? dirty_1_120 : _GEN_7382; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7931 = 3'h4 == state ? dirty_1_121 : _GEN_7383; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7932 = 3'h4 == state ? dirty_1_122 : _GEN_7384; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7933 = 3'h4 == state ? dirty_1_123 : _GEN_7385; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7934 = 3'h4 == state ? dirty_1_124 : _GEN_7386; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7935 = 3'h4 == state ? dirty_1_125 : _GEN_7387; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7936 = 3'h4 == state ? dirty_1_126 : _GEN_7388; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7937 = 3'h4 == state ? dirty_1_127 : _GEN_7389; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7938 = 3'h4 == state ? dirty_1_128 : _GEN_7390; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7939 = 3'h4 == state ? dirty_1_129 : _GEN_7391; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7940 = 3'h4 == state ? dirty_1_130 : _GEN_7392; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7941 = 3'h4 == state ? dirty_1_131 : _GEN_7393; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7942 = 3'h4 == state ? dirty_1_132 : _GEN_7394; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7943 = 3'h4 == state ? dirty_1_133 : _GEN_7395; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7944 = 3'h4 == state ? dirty_1_134 : _GEN_7396; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7945 = 3'h4 == state ? dirty_1_135 : _GEN_7397; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7946 = 3'h4 == state ? dirty_1_136 : _GEN_7398; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7947 = 3'h4 == state ? dirty_1_137 : _GEN_7399; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7948 = 3'h4 == state ? dirty_1_138 : _GEN_7400; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7949 = 3'h4 == state ? dirty_1_139 : _GEN_7401; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7950 = 3'h4 == state ? dirty_1_140 : _GEN_7402; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7951 = 3'h4 == state ? dirty_1_141 : _GEN_7403; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7952 = 3'h4 == state ? dirty_1_142 : _GEN_7404; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7953 = 3'h4 == state ? dirty_1_143 : _GEN_7405; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7954 = 3'h4 == state ? dirty_1_144 : _GEN_7406; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7955 = 3'h4 == state ? dirty_1_145 : _GEN_7407; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7956 = 3'h4 == state ? dirty_1_146 : _GEN_7408; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7957 = 3'h4 == state ? dirty_1_147 : _GEN_7409; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7958 = 3'h4 == state ? dirty_1_148 : _GEN_7410; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7959 = 3'h4 == state ? dirty_1_149 : _GEN_7411; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7960 = 3'h4 == state ? dirty_1_150 : _GEN_7412; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7961 = 3'h4 == state ? dirty_1_151 : _GEN_7413; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7962 = 3'h4 == state ? dirty_1_152 : _GEN_7414; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7963 = 3'h4 == state ? dirty_1_153 : _GEN_7415; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7964 = 3'h4 == state ? dirty_1_154 : _GEN_7416; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7965 = 3'h4 == state ? dirty_1_155 : _GEN_7417; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7966 = 3'h4 == state ? dirty_1_156 : _GEN_7418; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7967 = 3'h4 == state ? dirty_1_157 : _GEN_7419; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7968 = 3'h4 == state ? dirty_1_158 : _GEN_7420; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7969 = 3'h4 == state ? dirty_1_159 : _GEN_7421; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7970 = 3'h4 == state ? dirty_1_160 : _GEN_7422; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7971 = 3'h4 == state ? dirty_1_161 : _GEN_7423; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7972 = 3'h4 == state ? dirty_1_162 : _GEN_7424; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7973 = 3'h4 == state ? dirty_1_163 : _GEN_7425; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7974 = 3'h4 == state ? dirty_1_164 : _GEN_7426; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7975 = 3'h4 == state ? dirty_1_165 : _GEN_7427; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7976 = 3'h4 == state ? dirty_1_166 : _GEN_7428; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7977 = 3'h4 == state ? dirty_1_167 : _GEN_7429; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7978 = 3'h4 == state ? dirty_1_168 : _GEN_7430; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7979 = 3'h4 == state ? dirty_1_169 : _GEN_7431; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7980 = 3'h4 == state ? dirty_1_170 : _GEN_7432; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7981 = 3'h4 == state ? dirty_1_171 : _GEN_7433; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7982 = 3'h4 == state ? dirty_1_172 : _GEN_7434; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7983 = 3'h4 == state ? dirty_1_173 : _GEN_7435; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7984 = 3'h4 == state ? dirty_1_174 : _GEN_7436; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7985 = 3'h4 == state ? dirty_1_175 : _GEN_7437; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7986 = 3'h4 == state ? dirty_1_176 : _GEN_7438; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7987 = 3'h4 == state ? dirty_1_177 : _GEN_7439; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7988 = 3'h4 == state ? dirty_1_178 : _GEN_7440; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7989 = 3'h4 == state ? dirty_1_179 : _GEN_7441; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7990 = 3'h4 == state ? dirty_1_180 : _GEN_7442; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7991 = 3'h4 == state ? dirty_1_181 : _GEN_7443; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7992 = 3'h4 == state ? dirty_1_182 : _GEN_7444; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7993 = 3'h4 == state ? dirty_1_183 : _GEN_7445; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7994 = 3'h4 == state ? dirty_1_184 : _GEN_7446; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7995 = 3'h4 == state ? dirty_1_185 : _GEN_7447; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7996 = 3'h4 == state ? dirty_1_186 : _GEN_7448; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7997 = 3'h4 == state ? dirty_1_187 : _GEN_7449; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7998 = 3'h4 == state ? dirty_1_188 : _GEN_7450; // @[dcache.scala 183:18 113:28]
  wire  _GEN_7999 = 3'h4 == state ? dirty_1_189 : _GEN_7451; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8000 = 3'h4 == state ? dirty_1_190 : _GEN_7452; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8001 = 3'h4 == state ? dirty_1_191 : _GEN_7453; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8002 = 3'h4 == state ? dirty_1_192 : _GEN_7454; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8003 = 3'h4 == state ? dirty_1_193 : _GEN_7455; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8004 = 3'h4 == state ? dirty_1_194 : _GEN_7456; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8005 = 3'h4 == state ? dirty_1_195 : _GEN_7457; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8006 = 3'h4 == state ? dirty_1_196 : _GEN_7458; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8007 = 3'h4 == state ? dirty_1_197 : _GEN_7459; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8008 = 3'h4 == state ? dirty_1_198 : _GEN_7460; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8009 = 3'h4 == state ? dirty_1_199 : _GEN_7461; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8010 = 3'h4 == state ? dirty_1_200 : _GEN_7462; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8011 = 3'h4 == state ? dirty_1_201 : _GEN_7463; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8012 = 3'h4 == state ? dirty_1_202 : _GEN_7464; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8013 = 3'h4 == state ? dirty_1_203 : _GEN_7465; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8014 = 3'h4 == state ? dirty_1_204 : _GEN_7466; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8015 = 3'h4 == state ? dirty_1_205 : _GEN_7467; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8016 = 3'h4 == state ? dirty_1_206 : _GEN_7468; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8017 = 3'h4 == state ? dirty_1_207 : _GEN_7469; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8018 = 3'h4 == state ? dirty_1_208 : _GEN_7470; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8019 = 3'h4 == state ? dirty_1_209 : _GEN_7471; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8020 = 3'h4 == state ? dirty_1_210 : _GEN_7472; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8021 = 3'h4 == state ? dirty_1_211 : _GEN_7473; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8022 = 3'h4 == state ? dirty_1_212 : _GEN_7474; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8023 = 3'h4 == state ? dirty_1_213 : _GEN_7475; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8024 = 3'h4 == state ? dirty_1_214 : _GEN_7476; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8025 = 3'h4 == state ? dirty_1_215 : _GEN_7477; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8026 = 3'h4 == state ? dirty_1_216 : _GEN_7478; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8027 = 3'h4 == state ? dirty_1_217 : _GEN_7479; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8028 = 3'h4 == state ? dirty_1_218 : _GEN_7480; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8029 = 3'h4 == state ? dirty_1_219 : _GEN_7481; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8030 = 3'h4 == state ? dirty_1_220 : _GEN_7482; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8031 = 3'h4 == state ? dirty_1_221 : _GEN_7483; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8032 = 3'h4 == state ? dirty_1_222 : _GEN_7484; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8033 = 3'h4 == state ? dirty_1_223 : _GEN_7485; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8034 = 3'h4 == state ? dirty_1_224 : _GEN_7486; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8035 = 3'h4 == state ? dirty_1_225 : _GEN_7487; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8036 = 3'h4 == state ? dirty_1_226 : _GEN_7488; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8037 = 3'h4 == state ? dirty_1_227 : _GEN_7489; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8038 = 3'h4 == state ? dirty_1_228 : _GEN_7490; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8039 = 3'h4 == state ? dirty_1_229 : _GEN_7491; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8040 = 3'h4 == state ? dirty_1_230 : _GEN_7492; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8041 = 3'h4 == state ? dirty_1_231 : _GEN_7493; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8042 = 3'h4 == state ? dirty_1_232 : _GEN_7494; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8043 = 3'h4 == state ? dirty_1_233 : _GEN_7495; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8044 = 3'h4 == state ? dirty_1_234 : _GEN_7496; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8045 = 3'h4 == state ? dirty_1_235 : _GEN_7497; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8046 = 3'h4 == state ? dirty_1_236 : _GEN_7498; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8047 = 3'h4 == state ? dirty_1_237 : _GEN_7499; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8048 = 3'h4 == state ? dirty_1_238 : _GEN_7500; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8049 = 3'h4 == state ? dirty_1_239 : _GEN_7501; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8050 = 3'h4 == state ? dirty_1_240 : _GEN_7502; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8051 = 3'h4 == state ? dirty_1_241 : _GEN_7503; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8052 = 3'h4 == state ? dirty_1_242 : _GEN_7504; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8053 = 3'h4 == state ? dirty_1_243 : _GEN_7505; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8054 = 3'h4 == state ? dirty_1_244 : _GEN_7506; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8055 = 3'h4 == state ? dirty_1_245 : _GEN_7507; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8056 = 3'h4 == state ? dirty_1_246 : _GEN_7508; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8057 = 3'h4 == state ? dirty_1_247 : _GEN_7509; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8058 = 3'h4 == state ? dirty_1_248 : _GEN_7510; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8059 = 3'h4 == state ? dirty_1_249 : _GEN_7511; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8060 = 3'h4 == state ? dirty_1_250 : _GEN_7512; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8061 = 3'h4 == state ? dirty_1_251 : _GEN_7513; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8062 = 3'h4 == state ? dirty_1_252 : _GEN_7514; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8063 = 3'h4 == state ? dirty_1_253 : _GEN_7515; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8064 = 3'h4 == state ? dirty_1_254 : _GEN_7516; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8065 = 3'h4 == state ? dirty_1_255 : _GEN_7517; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8066 = 3'h4 == state ? 1'h0 : 3'h5 == state & _GEN_6973; // @[dcache.scala 183:18 144:25]
  wire  _GEN_8067 = 3'h4 == state ? 1'h0 : 3'h5 == state & _GEN_6974; // @[dcache.scala 183:18 144:25]
  wire [20:0] _GEN_8068 = 3'h4 == state ? 21'h0 : _GEN_7520; // @[dcache.scala 183:18 143:25]
  wire [20:0] _GEN_8069 = 3'h4 == state ? 21'h0 : _GEN_7521; // @[dcache.scala 183:18 143:25]
  wire  _GEN_8070 = 3'h4 == state ? 1'h0 : 3'h5 == state & _GEN_6977; // @[dcache.scala 183:18 157:25]
  wire [31:0] _GEN_8071 = 3'h4 == state ? 32'h7777 : _GEN_7523; // @[dcache.scala 183:18 155:25]
  wire  _GEN_8072 = 3'h4 == state ? req_valid : _GEN_7524; // @[dcache.scala 183:18 116:34]
  wire  _GEN_8073 = 3'h4 == state ? 1'h0 : 3'h5 == state & _GEN_6980; // @[dcache.scala 183:18 97:21]
  wire [21:0] _GEN_8074 = 3'h4 == state ? 22'h0 : _GEN_7526; // @[dcache.scala 183:18 98:21]
  wire  _GEN_8075 = 3'h4 == state ? cacheInst_r : _GEN_7527; // @[dcache.scala 183:18 89:38]
  wire  _GEN_8076 = 3'h4 == state ? invalidate : _GEN_7528; // @[dcache.scala 183:18 90:38]
  wire  _GEN_8077 = 3'h4 == state ? indexOnly : _GEN_7529; // @[dcache.scala 183:18 94:38]
  wire  _GEN_8078 = 3'h4 == state ? writeBack : _GEN_7530; // @[dcache.scala 183:18 93:38]
  wire  _GEN_8079 = 3'h4 == state ? storeTag : _GEN_7531; // @[dcache.scala 183:18 92:38]
  wire  _GEN_8080 = 3'h4 == state ? loadTag : _GEN_7532; // @[dcache.scala 183:18 91:38]
  wire [2:0] _GEN_8081 = 3'h3 == state ? _GEN_705 : _GEN_7533; // @[dcache.scala 183:18]
  wire [31:0] _GEN_8084 = 3'h3 == state ? _GEN_707 : 32'h0; // @[dcache.scala 183:18 163:25]
  wire [127:0] _GEN_8085 = 3'h3 == state ? _GEN_708 : 128'h0; // @[dcache.scala 183:18 165:25]
  wire [2:0] _GEN_8086 = 3'h3 == state ? _GEN_709 : 3'h0; // @[dcache.scala 183:18 162:25]
  wire [3:0] _GEN_8087 = 3'h3 == state ? _GEN_710 : 4'h0; // @[dcache.scala 183:18 164:25]
  wire  _GEN_8088 = 3'h3 == state ? _GEN_711 : _GEN_8070; // @[dcache.scala 183:18]
  wire  _GEN_8089 = 3'h3 == state ? 1'h0 : 3'h4 == state & _GEN_714; // @[dcache.scala 183:18 158:25]
  wire [2:0] _GEN_8090 = 3'h3 == state ? 3'h0 : _GEN_7535; // @[dcache.scala 183:18 159:25]
  wire [31:0] _GEN_8091 = 3'h3 == state ? 32'h0 : _GEN_7536; // @[dcache.scala 183:18 160:25]
  wire [1:0] _GEN_8092 = 3'h3 == state ? wr_cnt : _GEN_7537; // @[dcache.scala 183:18 178:34]
  wire [31:0] _GEN_8093 = 3'h3 == state ? 32'h0 : _GEN_7538; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8094 = 3'h3 == state ? 32'h0 : _GEN_7539; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8095 = 3'h3 == state ? 32'h0 : _GEN_7540; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8096 = 3'h3 == state ? 32'h0 : _GEN_7541; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8097 = 3'h3 == state ? 32'h0 : _GEN_7542; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8098 = 3'h3 == state ? 32'h0 : _GEN_7543; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8099 = 3'h3 == state ? 32'h0 : _GEN_7544; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8100 = 3'h3 == state ? 32'h0 : _GEN_7545; // @[dcache.scala 183:18 149:33]
  wire [3:0] _GEN_8101 = 3'h3 == state ? 4'h0 : _GEN_7546; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8102 = 3'h3 == state ? 4'h0 : _GEN_7547; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8103 = 3'h3 == state ? 4'h0 : _GEN_7548; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8104 = 3'h3 == state ? 4'h0 : _GEN_7549; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8105 = 3'h3 == state ? 4'h0 : _GEN_7550; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8106 = 3'h3 == state ? 4'h0 : _GEN_7551; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8107 = 3'h3 == state ? 4'h0 : _GEN_7552; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8108 = 3'h3 == state ? 4'h0 : _GEN_7553; // @[dcache.scala 183:18 150:33]
  wire  _GEN_8109 = 3'h3 == state ? dirty_0_0 : _GEN_7554; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8110 = 3'h3 == state ? dirty_0_1 : _GEN_7555; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8111 = 3'h3 == state ? dirty_0_2 : _GEN_7556; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8112 = 3'h3 == state ? dirty_0_3 : _GEN_7557; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8113 = 3'h3 == state ? dirty_0_4 : _GEN_7558; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8114 = 3'h3 == state ? dirty_0_5 : _GEN_7559; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8115 = 3'h3 == state ? dirty_0_6 : _GEN_7560; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8116 = 3'h3 == state ? dirty_0_7 : _GEN_7561; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8117 = 3'h3 == state ? dirty_0_8 : _GEN_7562; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8118 = 3'h3 == state ? dirty_0_9 : _GEN_7563; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8119 = 3'h3 == state ? dirty_0_10 : _GEN_7564; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8120 = 3'h3 == state ? dirty_0_11 : _GEN_7565; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8121 = 3'h3 == state ? dirty_0_12 : _GEN_7566; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8122 = 3'h3 == state ? dirty_0_13 : _GEN_7567; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8123 = 3'h3 == state ? dirty_0_14 : _GEN_7568; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8124 = 3'h3 == state ? dirty_0_15 : _GEN_7569; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8125 = 3'h3 == state ? dirty_0_16 : _GEN_7570; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8126 = 3'h3 == state ? dirty_0_17 : _GEN_7571; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8127 = 3'h3 == state ? dirty_0_18 : _GEN_7572; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8128 = 3'h3 == state ? dirty_0_19 : _GEN_7573; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8129 = 3'h3 == state ? dirty_0_20 : _GEN_7574; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8130 = 3'h3 == state ? dirty_0_21 : _GEN_7575; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8131 = 3'h3 == state ? dirty_0_22 : _GEN_7576; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8132 = 3'h3 == state ? dirty_0_23 : _GEN_7577; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8133 = 3'h3 == state ? dirty_0_24 : _GEN_7578; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8134 = 3'h3 == state ? dirty_0_25 : _GEN_7579; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8135 = 3'h3 == state ? dirty_0_26 : _GEN_7580; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8136 = 3'h3 == state ? dirty_0_27 : _GEN_7581; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8137 = 3'h3 == state ? dirty_0_28 : _GEN_7582; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8138 = 3'h3 == state ? dirty_0_29 : _GEN_7583; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8139 = 3'h3 == state ? dirty_0_30 : _GEN_7584; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8140 = 3'h3 == state ? dirty_0_31 : _GEN_7585; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8141 = 3'h3 == state ? dirty_0_32 : _GEN_7586; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8142 = 3'h3 == state ? dirty_0_33 : _GEN_7587; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8143 = 3'h3 == state ? dirty_0_34 : _GEN_7588; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8144 = 3'h3 == state ? dirty_0_35 : _GEN_7589; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8145 = 3'h3 == state ? dirty_0_36 : _GEN_7590; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8146 = 3'h3 == state ? dirty_0_37 : _GEN_7591; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8147 = 3'h3 == state ? dirty_0_38 : _GEN_7592; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8148 = 3'h3 == state ? dirty_0_39 : _GEN_7593; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8149 = 3'h3 == state ? dirty_0_40 : _GEN_7594; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8150 = 3'h3 == state ? dirty_0_41 : _GEN_7595; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8151 = 3'h3 == state ? dirty_0_42 : _GEN_7596; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8152 = 3'h3 == state ? dirty_0_43 : _GEN_7597; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8153 = 3'h3 == state ? dirty_0_44 : _GEN_7598; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8154 = 3'h3 == state ? dirty_0_45 : _GEN_7599; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8155 = 3'h3 == state ? dirty_0_46 : _GEN_7600; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8156 = 3'h3 == state ? dirty_0_47 : _GEN_7601; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8157 = 3'h3 == state ? dirty_0_48 : _GEN_7602; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8158 = 3'h3 == state ? dirty_0_49 : _GEN_7603; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8159 = 3'h3 == state ? dirty_0_50 : _GEN_7604; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8160 = 3'h3 == state ? dirty_0_51 : _GEN_7605; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8161 = 3'h3 == state ? dirty_0_52 : _GEN_7606; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8162 = 3'h3 == state ? dirty_0_53 : _GEN_7607; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8163 = 3'h3 == state ? dirty_0_54 : _GEN_7608; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8164 = 3'h3 == state ? dirty_0_55 : _GEN_7609; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8165 = 3'h3 == state ? dirty_0_56 : _GEN_7610; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8166 = 3'h3 == state ? dirty_0_57 : _GEN_7611; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8167 = 3'h3 == state ? dirty_0_58 : _GEN_7612; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8168 = 3'h3 == state ? dirty_0_59 : _GEN_7613; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8169 = 3'h3 == state ? dirty_0_60 : _GEN_7614; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8170 = 3'h3 == state ? dirty_0_61 : _GEN_7615; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8171 = 3'h3 == state ? dirty_0_62 : _GEN_7616; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8172 = 3'h3 == state ? dirty_0_63 : _GEN_7617; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8173 = 3'h3 == state ? dirty_0_64 : _GEN_7618; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8174 = 3'h3 == state ? dirty_0_65 : _GEN_7619; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8175 = 3'h3 == state ? dirty_0_66 : _GEN_7620; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8176 = 3'h3 == state ? dirty_0_67 : _GEN_7621; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8177 = 3'h3 == state ? dirty_0_68 : _GEN_7622; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8178 = 3'h3 == state ? dirty_0_69 : _GEN_7623; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8179 = 3'h3 == state ? dirty_0_70 : _GEN_7624; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8180 = 3'h3 == state ? dirty_0_71 : _GEN_7625; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8181 = 3'h3 == state ? dirty_0_72 : _GEN_7626; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8182 = 3'h3 == state ? dirty_0_73 : _GEN_7627; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8183 = 3'h3 == state ? dirty_0_74 : _GEN_7628; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8184 = 3'h3 == state ? dirty_0_75 : _GEN_7629; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8185 = 3'h3 == state ? dirty_0_76 : _GEN_7630; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8186 = 3'h3 == state ? dirty_0_77 : _GEN_7631; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8187 = 3'h3 == state ? dirty_0_78 : _GEN_7632; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8188 = 3'h3 == state ? dirty_0_79 : _GEN_7633; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8189 = 3'h3 == state ? dirty_0_80 : _GEN_7634; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8190 = 3'h3 == state ? dirty_0_81 : _GEN_7635; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8191 = 3'h3 == state ? dirty_0_82 : _GEN_7636; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8192 = 3'h3 == state ? dirty_0_83 : _GEN_7637; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8193 = 3'h3 == state ? dirty_0_84 : _GEN_7638; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8194 = 3'h3 == state ? dirty_0_85 : _GEN_7639; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8195 = 3'h3 == state ? dirty_0_86 : _GEN_7640; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8196 = 3'h3 == state ? dirty_0_87 : _GEN_7641; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8197 = 3'h3 == state ? dirty_0_88 : _GEN_7642; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8198 = 3'h3 == state ? dirty_0_89 : _GEN_7643; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8199 = 3'h3 == state ? dirty_0_90 : _GEN_7644; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8200 = 3'h3 == state ? dirty_0_91 : _GEN_7645; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8201 = 3'h3 == state ? dirty_0_92 : _GEN_7646; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8202 = 3'h3 == state ? dirty_0_93 : _GEN_7647; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8203 = 3'h3 == state ? dirty_0_94 : _GEN_7648; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8204 = 3'h3 == state ? dirty_0_95 : _GEN_7649; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8205 = 3'h3 == state ? dirty_0_96 : _GEN_7650; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8206 = 3'h3 == state ? dirty_0_97 : _GEN_7651; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8207 = 3'h3 == state ? dirty_0_98 : _GEN_7652; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8208 = 3'h3 == state ? dirty_0_99 : _GEN_7653; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8209 = 3'h3 == state ? dirty_0_100 : _GEN_7654; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8210 = 3'h3 == state ? dirty_0_101 : _GEN_7655; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8211 = 3'h3 == state ? dirty_0_102 : _GEN_7656; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8212 = 3'h3 == state ? dirty_0_103 : _GEN_7657; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8213 = 3'h3 == state ? dirty_0_104 : _GEN_7658; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8214 = 3'h3 == state ? dirty_0_105 : _GEN_7659; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8215 = 3'h3 == state ? dirty_0_106 : _GEN_7660; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8216 = 3'h3 == state ? dirty_0_107 : _GEN_7661; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8217 = 3'h3 == state ? dirty_0_108 : _GEN_7662; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8218 = 3'h3 == state ? dirty_0_109 : _GEN_7663; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8219 = 3'h3 == state ? dirty_0_110 : _GEN_7664; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8220 = 3'h3 == state ? dirty_0_111 : _GEN_7665; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8221 = 3'h3 == state ? dirty_0_112 : _GEN_7666; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8222 = 3'h3 == state ? dirty_0_113 : _GEN_7667; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8223 = 3'h3 == state ? dirty_0_114 : _GEN_7668; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8224 = 3'h3 == state ? dirty_0_115 : _GEN_7669; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8225 = 3'h3 == state ? dirty_0_116 : _GEN_7670; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8226 = 3'h3 == state ? dirty_0_117 : _GEN_7671; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8227 = 3'h3 == state ? dirty_0_118 : _GEN_7672; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8228 = 3'h3 == state ? dirty_0_119 : _GEN_7673; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8229 = 3'h3 == state ? dirty_0_120 : _GEN_7674; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8230 = 3'h3 == state ? dirty_0_121 : _GEN_7675; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8231 = 3'h3 == state ? dirty_0_122 : _GEN_7676; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8232 = 3'h3 == state ? dirty_0_123 : _GEN_7677; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8233 = 3'h3 == state ? dirty_0_124 : _GEN_7678; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8234 = 3'h3 == state ? dirty_0_125 : _GEN_7679; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8235 = 3'h3 == state ? dirty_0_126 : _GEN_7680; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8236 = 3'h3 == state ? dirty_0_127 : _GEN_7681; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8237 = 3'h3 == state ? dirty_0_128 : _GEN_7682; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8238 = 3'h3 == state ? dirty_0_129 : _GEN_7683; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8239 = 3'h3 == state ? dirty_0_130 : _GEN_7684; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8240 = 3'h3 == state ? dirty_0_131 : _GEN_7685; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8241 = 3'h3 == state ? dirty_0_132 : _GEN_7686; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8242 = 3'h3 == state ? dirty_0_133 : _GEN_7687; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8243 = 3'h3 == state ? dirty_0_134 : _GEN_7688; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8244 = 3'h3 == state ? dirty_0_135 : _GEN_7689; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8245 = 3'h3 == state ? dirty_0_136 : _GEN_7690; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8246 = 3'h3 == state ? dirty_0_137 : _GEN_7691; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8247 = 3'h3 == state ? dirty_0_138 : _GEN_7692; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8248 = 3'h3 == state ? dirty_0_139 : _GEN_7693; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8249 = 3'h3 == state ? dirty_0_140 : _GEN_7694; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8250 = 3'h3 == state ? dirty_0_141 : _GEN_7695; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8251 = 3'h3 == state ? dirty_0_142 : _GEN_7696; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8252 = 3'h3 == state ? dirty_0_143 : _GEN_7697; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8253 = 3'h3 == state ? dirty_0_144 : _GEN_7698; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8254 = 3'h3 == state ? dirty_0_145 : _GEN_7699; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8255 = 3'h3 == state ? dirty_0_146 : _GEN_7700; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8256 = 3'h3 == state ? dirty_0_147 : _GEN_7701; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8257 = 3'h3 == state ? dirty_0_148 : _GEN_7702; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8258 = 3'h3 == state ? dirty_0_149 : _GEN_7703; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8259 = 3'h3 == state ? dirty_0_150 : _GEN_7704; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8260 = 3'h3 == state ? dirty_0_151 : _GEN_7705; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8261 = 3'h3 == state ? dirty_0_152 : _GEN_7706; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8262 = 3'h3 == state ? dirty_0_153 : _GEN_7707; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8263 = 3'h3 == state ? dirty_0_154 : _GEN_7708; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8264 = 3'h3 == state ? dirty_0_155 : _GEN_7709; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8265 = 3'h3 == state ? dirty_0_156 : _GEN_7710; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8266 = 3'h3 == state ? dirty_0_157 : _GEN_7711; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8267 = 3'h3 == state ? dirty_0_158 : _GEN_7712; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8268 = 3'h3 == state ? dirty_0_159 : _GEN_7713; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8269 = 3'h3 == state ? dirty_0_160 : _GEN_7714; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8270 = 3'h3 == state ? dirty_0_161 : _GEN_7715; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8271 = 3'h3 == state ? dirty_0_162 : _GEN_7716; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8272 = 3'h3 == state ? dirty_0_163 : _GEN_7717; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8273 = 3'h3 == state ? dirty_0_164 : _GEN_7718; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8274 = 3'h3 == state ? dirty_0_165 : _GEN_7719; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8275 = 3'h3 == state ? dirty_0_166 : _GEN_7720; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8276 = 3'h3 == state ? dirty_0_167 : _GEN_7721; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8277 = 3'h3 == state ? dirty_0_168 : _GEN_7722; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8278 = 3'h3 == state ? dirty_0_169 : _GEN_7723; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8279 = 3'h3 == state ? dirty_0_170 : _GEN_7724; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8280 = 3'h3 == state ? dirty_0_171 : _GEN_7725; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8281 = 3'h3 == state ? dirty_0_172 : _GEN_7726; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8282 = 3'h3 == state ? dirty_0_173 : _GEN_7727; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8283 = 3'h3 == state ? dirty_0_174 : _GEN_7728; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8284 = 3'h3 == state ? dirty_0_175 : _GEN_7729; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8285 = 3'h3 == state ? dirty_0_176 : _GEN_7730; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8286 = 3'h3 == state ? dirty_0_177 : _GEN_7731; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8287 = 3'h3 == state ? dirty_0_178 : _GEN_7732; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8288 = 3'h3 == state ? dirty_0_179 : _GEN_7733; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8289 = 3'h3 == state ? dirty_0_180 : _GEN_7734; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8290 = 3'h3 == state ? dirty_0_181 : _GEN_7735; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8291 = 3'h3 == state ? dirty_0_182 : _GEN_7736; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8292 = 3'h3 == state ? dirty_0_183 : _GEN_7737; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8293 = 3'h3 == state ? dirty_0_184 : _GEN_7738; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8294 = 3'h3 == state ? dirty_0_185 : _GEN_7739; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8295 = 3'h3 == state ? dirty_0_186 : _GEN_7740; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8296 = 3'h3 == state ? dirty_0_187 : _GEN_7741; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8297 = 3'h3 == state ? dirty_0_188 : _GEN_7742; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8298 = 3'h3 == state ? dirty_0_189 : _GEN_7743; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8299 = 3'h3 == state ? dirty_0_190 : _GEN_7744; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8300 = 3'h3 == state ? dirty_0_191 : _GEN_7745; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8301 = 3'h3 == state ? dirty_0_192 : _GEN_7746; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8302 = 3'h3 == state ? dirty_0_193 : _GEN_7747; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8303 = 3'h3 == state ? dirty_0_194 : _GEN_7748; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8304 = 3'h3 == state ? dirty_0_195 : _GEN_7749; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8305 = 3'h3 == state ? dirty_0_196 : _GEN_7750; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8306 = 3'h3 == state ? dirty_0_197 : _GEN_7751; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8307 = 3'h3 == state ? dirty_0_198 : _GEN_7752; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8308 = 3'h3 == state ? dirty_0_199 : _GEN_7753; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8309 = 3'h3 == state ? dirty_0_200 : _GEN_7754; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8310 = 3'h3 == state ? dirty_0_201 : _GEN_7755; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8311 = 3'h3 == state ? dirty_0_202 : _GEN_7756; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8312 = 3'h3 == state ? dirty_0_203 : _GEN_7757; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8313 = 3'h3 == state ? dirty_0_204 : _GEN_7758; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8314 = 3'h3 == state ? dirty_0_205 : _GEN_7759; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8315 = 3'h3 == state ? dirty_0_206 : _GEN_7760; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8316 = 3'h3 == state ? dirty_0_207 : _GEN_7761; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8317 = 3'h3 == state ? dirty_0_208 : _GEN_7762; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8318 = 3'h3 == state ? dirty_0_209 : _GEN_7763; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8319 = 3'h3 == state ? dirty_0_210 : _GEN_7764; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8320 = 3'h3 == state ? dirty_0_211 : _GEN_7765; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8321 = 3'h3 == state ? dirty_0_212 : _GEN_7766; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8322 = 3'h3 == state ? dirty_0_213 : _GEN_7767; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8323 = 3'h3 == state ? dirty_0_214 : _GEN_7768; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8324 = 3'h3 == state ? dirty_0_215 : _GEN_7769; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8325 = 3'h3 == state ? dirty_0_216 : _GEN_7770; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8326 = 3'h3 == state ? dirty_0_217 : _GEN_7771; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8327 = 3'h3 == state ? dirty_0_218 : _GEN_7772; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8328 = 3'h3 == state ? dirty_0_219 : _GEN_7773; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8329 = 3'h3 == state ? dirty_0_220 : _GEN_7774; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8330 = 3'h3 == state ? dirty_0_221 : _GEN_7775; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8331 = 3'h3 == state ? dirty_0_222 : _GEN_7776; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8332 = 3'h3 == state ? dirty_0_223 : _GEN_7777; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8333 = 3'h3 == state ? dirty_0_224 : _GEN_7778; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8334 = 3'h3 == state ? dirty_0_225 : _GEN_7779; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8335 = 3'h3 == state ? dirty_0_226 : _GEN_7780; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8336 = 3'h3 == state ? dirty_0_227 : _GEN_7781; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8337 = 3'h3 == state ? dirty_0_228 : _GEN_7782; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8338 = 3'h3 == state ? dirty_0_229 : _GEN_7783; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8339 = 3'h3 == state ? dirty_0_230 : _GEN_7784; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8340 = 3'h3 == state ? dirty_0_231 : _GEN_7785; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8341 = 3'h3 == state ? dirty_0_232 : _GEN_7786; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8342 = 3'h3 == state ? dirty_0_233 : _GEN_7787; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8343 = 3'h3 == state ? dirty_0_234 : _GEN_7788; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8344 = 3'h3 == state ? dirty_0_235 : _GEN_7789; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8345 = 3'h3 == state ? dirty_0_236 : _GEN_7790; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8346 = 3'h3 == state ? dirty_0_237 : _GEN_7791; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8347 = 3'h3 == state ? dirty_0_238 : _GEN_7792; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8348 = 3'h3 == state ? dirty_0_239 : _GEN_7793; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8349 = 3'h3 == state ? dirty_0_240 : _GEN_7794; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8350 = 3'h3 == state ? dirty_0_241 : _GEN_7795; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8351 = 3'h3 == state ? dirty_0_242 : _GEN_7796; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8352 = 3'h3 == state ? dirty_0_243 : _GEN_7797; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8353 = 3'h3 == state ? dirty_0_244 : _GEN_7798; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8354 = 3'h3 == state ? dirty_0_245 : _GEN_7799; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8355 = 3'h3 == state ? dirty_0_246 : _GEN_7800; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8356 = 3'h3 == state ? dirty_0_247 : _GEN_7801; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8357 = 3'h3 == state ? dirty_0_248 : _GEN_7802; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8358 = 3'h3 == state ? dirty_0_249 : _GEN_7803; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8359 = 3'h3 == state ? dirty_0_250 : _GEN_7804; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8360 = 3'h3 == state ? dirty_0_251 : _GEN_7805; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8361 = 3'h3 == state ? dirty_0_252 : _GEN_7806; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8362 = 3'h3 == state ? dirty_0_253 : _GEN_7807; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8363 = 3'h3 == state ? dirty_0_254 : _GEN_7808; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8364 = 3'h3 == state ? dirty_0_255 : _GEN_7809; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8365 = 3'h3 == state ? dirty_1_0 : _GEN_7810; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8366 = 3'h3 == state ? dirty_1_1 : _GEN_7811; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8367 = 3'h3 == state ? dirty_1_2 : _GEN_7812; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8368 = 3'h3 == state ? dirty_1_3 : _GEN_7813; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8369 = 3'h3 == state ? dirty_1_4 : _GEN_7814; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8370 = 3'h3 == state ? dirty_1_5 : _GEN_7815; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8371 = 3'h3 == state ? dirty_1_6 : _GEN_7816; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8372 = 3'h3 == state ? dirty_1_7 : _GEN_7817; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8373 = 3'h3 == state ? dirty_1_8 : _GEN_7818; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8374 = 3'h3 == state ? dirty_1_9 : _GEN_7819; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8375 = 3'h3 == state ? dirty_1_10 : _GEN_7820; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8376 = 3'h3 == state ? dirty_1_11 : _GEN_7821; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8377 = 3'h3 == state ? dirty_1_12 : _GEN_7822; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8378 = 3'h3 == state ? dirty_1_13 : _GEN_7823; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8379 = 3'h3 == state ? dirty_1_14 : _GEN_7824; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8380 = 3'h3 == state ? dirty_1_15 : _GEN_7825; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8381 = 3'h3 == state ? dirty_1_16 : _GEN_7826; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8382 = 3'h3 == state ? dirty_1_17 : _GEN_7827; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8383 = 3'h3 == state ? dirty_1_18 : _GEN_7828; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8384 = 3'h3 == state ? dirty_1_19 : _GEN_7829; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8385 = 3'h3 == state ? dirty_1_20 : _GEN_7830; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8386 = 3'h3 == state ? dirty_1_21 : _GEN_7831; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8387 = 3'h3 == state ? dirty_1_22 : _GEN_7832; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8388 = 3'h3 == state ? dirty_1_23 : _GEN_7833; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8389 = 3'h3 == state ? dirty_1_24 : _GEN_7834; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8390 = 3'h3 == state ? dirty_1_25 : _GEN_7835; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8391 = 3'h3 == state ? dirty_1_26 : _GEN_7836; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8392 = 3'h3 == state ? dirty_1_27 : _GEN_7837; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8393 = 3'h3 == state ? dirty_1_28 : _GEN_7838; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8394 = 3'h3 == state ? dirty_1_29 : _GEN_7839; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8395 = 3'h3 == state ? dirty_1_30 : _GEN_7840; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8396 = 3'h3 == state ? dirty_1_31 : _GEN_7841; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8397 = 3'h3 == state ? dirty_1_32 : _GEN_7842; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8398 = 3'h3 == state ? dirty_1_33 : _GEN_7843; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8399 = 3'h3 == state ? dirty_1_34 : _GEN_7844; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8400 = 3'h3 == state ? dirty_1_35 : _GEN_7845; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8401 = 3'h3 == state ? dirty_1_36 : _GEN_7846; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8402 = 3'h3 == state ? dirty_1_37 : _GEN_7847; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8403 = 3'h3 == state ? dirty_1_38 : _GEN_7848; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8404 = 3'h3 == state ? dirty_1_39 : _GEN_7849; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8405 = 3'h3 == state ? dirty_1_40 : _GEN_7850; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8406 = 3'h3 == state ? dirty_1_41 : _GEN_7851; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8407 = 3'h3 == state ? dirty_1_42 : _GEN_7852; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8408 = 3'h3 == state ? dirty_1_43 : _GEN_7853; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8409 = 3'h3 == state ? dirty_1_44 : _GEN_7854; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8410 = 3'h3 == state ? dirty_1_45 : _GEN_7855; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8411 = 3'h3 == state ? dirty_1_46 : _GEN_7856; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8412 = 3'h3 == state ? dirty_1_47 : _GEN_7857; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8413 = 3'h3 == state ? dirty_1_48 : _GEN_7858; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8414 = 3'h3 == state ? dirty_1_49 : _GEN_7859; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8415 = 3'h3 == state ? dirty_1_50 : _GEN_7860; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8416 = 3'h3 == state ? dirty_1_51 : _GEN_7861; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8417 = 3'h3 == state ? dirty_1_52 : _GEN_7862; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8418 = 3'h3 == state ? dirty_1_53 : _GEN_7863; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8419 = 3'h3 == state ? dirty_1_54 : _GEN_7864; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8420 = 3'h3 == state ? dirty_1_55 : _GEN_7865; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8421 = 3'h3 == state ? dirty_1_56 : _GEN_7866; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8422 = 3'h3 == state ? dirty_1_57 : _GEN_7867; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8423 = 3'h3 == state ? dirty_1_58 : _GEN_7868; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8424 = 3'h3 == state ? dirty_1_59 : _GEN_7869; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8425 = 3'h3 == state ? dirty_1_60 : _GEN_7870; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8426 = 3'h3 == state ? dirty_1_61 : _GEN_7871; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8427 = 3'h3 == state ? dirty_1_62 : _GEN_7872; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8428 = 3'h3 == state ? dirty_1_63 : _GEN_7873; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8429 = 3'h3 == state ? dirty_1_64 : _GEN_7874; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8430 = 3'h3 == state ? dirty_1_65 : _GEN_7875; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8431 = 3'h3 == state ? dirty_1_66 : _GEN_7876; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8432 = 3'h3 == state ? dirty_1_67 : _GEN_7877; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8433 = 3'h3 == state ? dirty_1_68 : _GEN_7878; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8434 = 3'h3 == state ? dirty_1_69 : _GEN_7879; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8435 = 3'h3 == state ? dirty_1_70 : _GEN_7880; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8436 = 3'h3 == state ? dirty_1_71 : _GEN_7881; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8437 = 3'h3 == state ? dirty_1_72 : _GEN_7882; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8438 = 3'h3 == state ? dirty_1_73 : _GEN_7883; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8439 = 3'h3 == state ? dirty_1_74 : _GEN_7884; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8440 = 3'h3 == state ? dirty_1_75 : _GEN_7885; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8441 = 3'h3 == state ? dirty_1_76 : _GEN_7886; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8442 = 3'h3 == state ? dirty_1_77 : _GEN_7887; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8443 = 3'h3 == state ? dirty_1_78 : _GEN_7888; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8444 = 3'h3 == state ? dirty_1_79 : _GEN_7889; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8445 = 3'h3 == state ? dirty_1_80 : _GEN_7890; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8446 = 3'h3 == state ? dirty_1_81 : _GEN_7891; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8447 = 3'h3 == state ? dirty_1_82 : _GEN_7892; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8448 = 3'h3 == state ? dirty_1_83 : _GEN_7893; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8449 = 3'h3 == state ? dirty_1_84 : _GEN_7894; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8450 = 3'h3 == state ? dirty_1_85 : _GEN_7895; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8451 = 3'h3 == state ? dirty_1_86 : _GEN_7896; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8452 = 3'h3 == state ? dirty_1_87 : _GEN_7897; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8453 = 3'h3 == state ? dirty_1_88 : _GEN_7898; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8454 = 3'h3 == state ? dirty_1_89 : _GEN_7899; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8455 = 3'h3 == state ? dirty_1_90 : _GEN_7900; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8456 = 3'h3 == state ? dirty_1_91 : _GEN_7901; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8457 = 3'h3 == state ? dirty_1_92 : _GEN_7902; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8458 = 3'h3 == state ? dirty_1_93 : _GEN_7903; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8459 = 3'h3 == state ? dirty_1_94 : _GEN_7904; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8460 = 3'h3 == state ? dirty_1_95 : _GEN_7905; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8461 = 3'h3 == state ? dirty_1_96 : _GEN_7906; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8462 = 3'h3 == state ? dirty_1_97 : _GEN_7907; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8463 = 3'h3 == state ? dirty_1_98 : _GEN_7908; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8464 = 3'h3 == state ? dirty_1_99 : _GEN_7909; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8465 = 3'h3 == state ? dirty_1_100 : _GEN_7910; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8466 = 3'h3 == state ? dirty_1_101 : _GEN_7911; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8467 = 3'h3 == state ? dirty_1_102 : _GEN_7912; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8468 = 3'h3 == state ? dirty_1_103 : _GEN_7913; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8469 = 3'h3 == state ? dirty_1_104 : _GEN_7914; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8470 = 3'h3 == state ? dirty_1_105 : _GEN_7915; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8471 = 3'h3 == state ? dirty_1_106 : _GEN_7916; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8472 = 3'h3 == state ? dirty_1_107 : _GEN_7917; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8473 = 3'h3 == state ? dirty_1_108 : _GEN_7918; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8474 = 3'h3 == state ? dirty_1_109 : _GEN_7919; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8475 = 3'h3 == state ? dirty_1_110 : _GEN_7920; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8476 = 3'h3 == state ? dirty_1_111 : _GEN_7921; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8477 = 3'h3 == state ? dirty_1_112 : _GEN_7922; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8478 = 3'h3 == state ? dirty_1_113 : _GEN_7923; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8479 = 3'h3 == state ? dirty_1_114 : _GEN_7924; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8480 = 3'h3 == state ? dirty_1_115 : _GEN_7925; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8481 = 3'h3 == state ? dirty_1_116 : _GEN_7926; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8482 = 3'h3 == state ? dirty_1_117 : _GEN_7927; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8483 = 3'h3 == state ? dirty_1_118 : _GEN_7928; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8484 = 3'h3 == state ? dirty_1_119 : _GEN_7929; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8485 = 3'h3 == state ? dirty_1_120 : _GEN_7930; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8486 = 3'h3 == state ? dirty_1_121 : _GEN_7931; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8487 = 3'h3 == state ? dirty_1_122 : _GEN_7932; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8488 = 3'h3 == state ? dirty_1_123 : _GEN_7933; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8489 = 3'h3 == state ? dirty_1_124 : _GEN_7934; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8490 = 3'h3 == state ? dirty_1_125 : _GEN_7935; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8491 = 3'h3 == state ? dirty_1_126 : _GEN_7936; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8492 = 3'h3 == state ? dirty_1_127 : _GEN_7937; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8493 = 3'h3 == state ? dirty_1_128 : _GEN_7938; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8494 = 3'h3 == state ? dirty_1_129 : _GEN_7939; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8495 = 3'h3 == state ? dirty_1_130 : _GEN_7940; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8496 = 3'h3 == state ? dirty_1_131 : _GEN_7941; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8497 = 3'h3 == state ? dirty_1_132 : _GEN_7942; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8498 = 3'h3 == state ? dirty_1_133 : _GEN_7943; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8499 = 3'h3 == state ? dirty_1_134 : _GEN_7944; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8500 = 3'h3 == state ? dirty_1_135 : _GEN_7945; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8501 = 3'h3 == state ? dirty_1_136 : _GEN_7946; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8502 = 3'h3 == state ? dirty_1_137 : _GEN_7947; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8503 = 3'h3 == state ? dirty_1_138 : _GEN_7948; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8504 = 3'h3 == state ? dirty_1_139 : _GEN_7949; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8505 = 3'h3 == state ? dirty_1_140 : _GEN_7950; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8506 = 3'h3 == state ? dirty_1_141 : _GEN_7951; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8507 = 3'h3 == state ? dirty_1_142 : _GEN_7952; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8508 = 3'h3 == state ? dirty_1_143 : _GEN_7953; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8509 = 3'h3 == state ? dirty_1_144 : _GEN_7954; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8510 = 3'h3 == state ? dirty_1_145 : _GEN_7955; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8511 = 3'h3 == state ? dirty_1_146 : _GEN_7956; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8512 = 3'h3 == state ? dirty_1_147 : _GEN_7957; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8513 = 3'h3 == state ? dirty_1_148 : _GEN_7958; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8514 = 3'h3 == state ? dirty_1_149 : _GEN_7959; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8515 = 3'h3 == state ? dirty_1_150 : _GEN_7960; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8516 = 3'h3 == state ? dirty_1_151 : _GEN_7961; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8517 = 3'h3 == state ? dirty_1_152 : _GEN_7962; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8518 = 3'h3 == state ? dirty_1_153 : _GEN_7963; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8519 = 3'h3 == state ? dirty_1_154 : _GEN_7964; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8520 = 3'h3 == state ? dirty_1_155 : _GEN_7965; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8521 = 3'h3 == state ? dirty_1_156 : _GEN_7966; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8522 = 3'h3 == state ? dirty_1_157 : _GEN_7967; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8523 = 3'h3 == state ? dirty_1_158 : _GEN_7968; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8524 = 3'h3 == state ? dirty_1_159 : _GEN_7969; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8525 = 3'h3 == state ? dirty_1_160 : _GEN_7970; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8526 = 3'h3 == state ? dirty_1_161 : _GEN_7971; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8527 = 3'h3 == state ? dirty_1_162 : _GEN_7972; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8528 = 3'h3 == state ? dirty_1_163 : _GEN_7973; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8529 = 3'h3 == state ? dirty_1_164 : _GEN_7974; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8530 = 3'h3 == state ? dirty_1_165 : _GEN_7975; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8531 = 3'h3 == state ? dirty_1_166 : _GEN_7976; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8532 = 3'h3 == state ? dirty_1_167 : _GEN_7977; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8533 = 3'h3 == state ? dirty_1_168 : _GEN_7978; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8534 = 3'h3 == state ? dirty_1_169 : _GEN_7979; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8535 = 3'h3 == state ? dirty_1_170 : _GEN_7980; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8536 = 3'h3 == state ? dirty_1_171 : _GEN_7981; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8537 = 3'h3 == state ? dirty_1_172 : _GEN_7982; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8538 = 3'h3 == state ? dirty_1_173 : _GEN_7983; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8539 = 3'h3 == state ? dirty_1_174 : _GEN_7984; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8540 = 3'h3 == state ? dirty_1_175 : _GEN_7985; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8541 = 3'h3 == state ? dirty_1_176 : _GEN_7986; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8542 = 3'h3 == state ? dirty_1_177 : _GEN_7987; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8543 = 3'h3 == state ? dirty_1_178 : _GEN_7988; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8544 = 3'h3 == state ? dirty_1_179 : _GEN_7989; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8545 = 3'h3 == state ? dirty_1_180 : _GEN_7990; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8546 = 3'h3 == state ? dirty_1_181 : _GEN_7991; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8547 = 3'h3 == state ? dirty_1_182 : _GEN_7992; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8548 = 3'h3 == state ? dirty_1_183 : _GEN_7993; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8549 = 3'h3 == state ? dirty_1_184 : _GEN_7994; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8550 = 3'h3 == state ? dirty_1_185 : _GEN_7995; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8551 = 3'h3 == state ? dirty_1_186 : _GEN_7996; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8552 = 3'h3 == state ? dirty_1_187 : _GEN_7997; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8553 = 3'h3 == state ? dirty_1_188 : _GEN_7998; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8554 = 3'h3 == state ? dirty_1_189 : _GEN_7999; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8555 = 3'h3 == state ? dirty_1_190 : _GEN_8000; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8556 = 3'h3 == state ? dirty_1_191 : _GEN_8001; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8557 = 3'h3 == state ? dirty_1_192 : _GEN_8002; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8558 = 3'h3 == state ? dirty_1_193 : _GEN_8003; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8559 = 3'h3 == state ? dirty_1_194 : _GEN_8004; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8560 = 3'h3 == state ? dirty_1_195 : _GEN_8005; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8561 = 3'h3 == state ? dirty_1_196 : _GEN_8006; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8562 = 3'h3 == state ? dirty_1_197 : _GEN_8007; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8563 = 3'h3 == state ? dirty_1_198 : _GEN_8008; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8564 = 3'h3 == state ? dirty_1_199 : _GEN_8009; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8565 = 3'h3 == state ? dirty_1_200 : _GEN_8010; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8566 = 3'h3 == state ? dirty_1_201 : _GEN_8011; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8567 = 3'h3 == state ? dirty_1_202 : _GEN_8012; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8568 = 3'h3 == state ? dirty_1_203 : _GEN_8013; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8569 = 3'h3 == state ? dirty_1_204 : _GEN_8014; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8570 = 3'h3 == state ? dirty_1_205 : _GEN_8015; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8571 = 3'h3 == state ? dirty_1_206 : _GEN_8016; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8572 = 3'h3 == state ? dirty_1_207 : _GEN_8017; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8573 = 3'h3 == state ? dirty_1_208 : _GEN_8018; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8574 = 3'h3 == state ? dirty_1_209 : _GEN_8019; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8575 = 3'h3 == state ? dirty_1_210 : _GEN_8020; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8576 = 3'h3 == state ? dirty_1_211 : _GEN_8021; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8577 = 3'h3 == state ? dirty_1_212 : _GEN_8022; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8578 = 3'h3 == state ? dirty_1_213 : _GEN_8023; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8579 = 3'h3 == state ? dirty_1_214 : _GEN_8024; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8580 = 3'h3 == state ? dirty_1_215 : _GEN_8025; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8581 = 3'h3 == state ? dirty_1_216 : _GEN_8026; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8582 = 3'h3 == state ? dirty_1_217 : _GEN_8027; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8583 = 3'h3 == state ? dirty_1_218 : _GEN_8028; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8584 = 3'h3 == state ? dirty_1_219 : _GEN_8029; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8585 = 3'h3 == state ? dirty_1_220 : _GEN_8030; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8586 = 3'h3 == state ? dirty_1_221 : _GEN_8031; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8587 = 3'h3 == state ? dirty_1_222 : _GEN_8032; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8588 = 3'h3 == state ? dirty_1_223 : _GEN_8033; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8589 = 3'h3 == state ? dirty_1_224 : _GEN_8034; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8590 = 3'h3 == state ? dirty_1_225 : _GEN_8035; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8591 = 3'h3 == state ? dirty_1_226 : _GEN_8036; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8592 = 3'h3 == state ? dirty_1_227 : _GEN_8037; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8593 = 3'h3 == state ? dirty_1_228 : _GEN_8038; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8594 = 3'h3 == state ? dirty_1_229 : _GEN_8039; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8595 = 3'h3 == state ? dirty_1_230 : _GEN_8040; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8596 = 3'h3 == state ? dirty_1_231 : _GEN_8041; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8597 = 3'h3 == state ? dirty_1_232 : _GEN_8042; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8598 = 3'h3 == state ? dirty_1_233 : _GEN_8043; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8599 = 3'h3 == state ? dirty_1_234 : _GEN_8044; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8600 = 3'h3 == state ? dirty_1_235 : _GEN_8045; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8601 = 3'h3 == state ? dirty_1_236 : _GEN_8046; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8602 = 3'h3 == state ? dirty_1_237 : _GEN_8047; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8603 = 3'h3 == state ? dirty_1_238 : _GEN_8048; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8604 = 3'h3 == state ? dirty_1_239 : _GEN_8049; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8605 = 3'h3 == state ? dirty_1_240 : _GEN_8050; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8606 = 3'h3 == state ? dirty_1_241 : _GEN_8051; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8607 = 3'h3 == state ? dirty_1_242 : _GEN_8052; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8608 = 3'h3 == state ? dirty_1_243 : _GEN_8053; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8609 = 3'h3 == state ? dirty_1_244 : _GEN_8054; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8610 = 3'h3 == state ? dirty_1_245 : _GEN_8055; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8611 = 3'h3 == state ? dirty_1_246 : _GEN_8056; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8612 = 3'h3 == state ? dirty_1_247 : _GEN_8057; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8613 = 3'h3 == state ? dirty_1_248 : _GEN_8058; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8614 = 3'h3 == state ? dirty_1_249 : _GEN_8059; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8615 = 3'h3 == state ? dirty_1_250 : _GEN_8060; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8616 = 3'h3 == state ? dirty_1_251 : _GEN_8061; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8617 = 3'h3 == state ? dirty_1_252 : _GEN_8062; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8618 = 3'h3 == state ? dirty_1_253 : _GEN_8063; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8619 = 3'h3 == state ? dirty_1_254 : _GEN_8064; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8620 = 3'h3 == state ? dirty_1_255 : _GEN_8065; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8621 = 3'h3 == state ? 1'h0 : _GEN_8066; // @[dcache.scala 183:18 144:25]
  wire  _GEN_8622 = 3'h3 == state ? 1'h0 : _GEN_8067; // @[dcache.scala 183:18 144:25]
  wire [20:0] _GEN_8623 = 3'h3 == state ? 21'h0 : _GEN_8068; // @[dcache.scala 183:18 143:25]
  wire [20:0] _GEN_8624 = 3'h3 == state ? 21'h0 : _GEN_8069; // @[dcache.scala 183:18 143:25]
  wire [31:0] _GEN_8625 = 3'h3 == state ? 32'h7777 : _GEN_8071; // @[dcache.scala 183:18 155:25]
  wire  _GEN_8626 = 3'h3 == state ? req_valid : _GEN_8072; // @[dcache.scala 183:18 116:34]
  wire  _GEN_8627 = 3'h3 == state ? 1'h0 : _GEN_8073; // @[dcache.scala 183:18 97:21]
  wire [21:0] _GEN_8628 = 3'h3 == state ? 22'h0 : _GEN_8074; // @[dcache.scala 183:18 98:21]
  wire  _GEN_8629 = 3'h3 == state ? cacheInst_r : _GEN_8075; // @[dcache.scala 183:18 89:38]
  wire  _GEN_8630 = 3'h3 == state ? invalidate : _GEN_8076; // @[dcache.scala 183:18 90:38]
  wire  _GEN_8631 = 3'h3 == state ? indexOnly : _GEN_8077; // @[dcache.scala 183:18 94:38]
  wire  _GEN_8632 = 3'h3 == state ? writeBack : _GEN_8078; // @[dcache.scala 183:18 93:38]
  wire  _GEN_8633 = 3'h3 == state ? storeTag : _GEN_8079; // @[dcache.scala 183:18 92:38]
  wire  _GEN_8634 = 3'h3 == state ? loadTag : _GEN_8080; // @[dcache.scala 183:18 91:38]
  wire  _GEN_9223 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_150; // @[dcache.scala 183:18 181:25]
  wire  refillIDX = 3'h0 == state ? 1'h0 : _GEN_9223; // @[dcache.scala 183:18 181:25]
  wire  _GEN_8640 = 3'h2 == state ? 1'h0 : 3'h3 == state & _GEN_706; // @[dcache.scala 183:18 161:25]
  wire [31:0] _GEN_8641 = 3'h2 == state ? 32'h0 : _GEN_8084; // @[dcache.scala 183:18 163:25]
  wire [127:0] _GEN_8642 = 3'h2 == state ? 128'h0 : _GEN_8085; // @[dcache.scala 183:18 165:25]
  wire [2:0] _GEN_8643 = 3'h2 == state ? 3'h0 : _GEN_8086; // @[dcache.scala 183:18 162:25]
  wire [3:0] _GEN_8644 = 3'h2 == state ? 4'h0 : _GEN_8087; // @[dcache.scala 183:18 164:25]
  wire  _GEN_8645 = 3'h2 == state ? 1'h0 : _GEN_8088; // @[dcache.scala 183:18 157:25]
  wire  _GEN_8646 = 3'h2 == state ? 1'h0 : _GEN_8089; // @[dcache.scala 183:18 158:25]
  wire [2:0] _GEN_8647 = 3'h2 == state ? 3'h0 : _GEN_8090; // @[dcache.scala 183:18 159:25]
  wire [31:0] _GEN_8648 = 3'h2 == state ? 32'h0 : _GEN_8091; // @[dcache.scala 183:18 160:25]
  wire [31:0] _GEN_8650 = 3'h2 == state ? 32'h0 : _GEN_8093; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8651 = 3'h2 == state ? 32'h0 : _GEN_8094; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8652 = 3'h2 == state ? 32'h0 : _GEN_8095; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8653 = 3'h2 == state ? 32'h0 : _GEN_8096; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8654 = 3'h2 == state ? 32'h0 : _GEN_8097; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8655 = 3'h2 == state ? 32'h0 : _GEN_8098; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8656 = 3'h2 == state ? 32'h0 : _GEN_8099; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_8657 = 3'h2 == state ? 32'h0 : _GEN_8100; // @[dcache.scala 183:18 149:33]
  wire [3:0] _GEN_8658 = 3'h2 == state ? 4'h0 : _GEN_8101; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8659 = 3'h2 == state ? 4'h0 : _GEN_8102; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8660 = 3'h2 == state ? 4'h0 : _GEN_8103; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8661 = 3'h2 == state ? 4'h0 : _GEN_8104; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8662 = 3'h2 == state ? 4'h0 : _GEN_8105; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8663 = 3'h2 == state ? 4'h0 : _GEN_8106; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8664 = 3'h2 == state ? 4'h0 : _GEN_8107; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_8665 = 3'h2 == state ? 4'h0 : _GEN_8108; // @[dcache.scala 183:18 150:33]
  wire  _GEN_8666 = 3'h2 == state ? dirty_0_0 : _GEN_8109; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8667 = 3'h2 == state ? dirty_0_1 : _GEN_8110; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8668 = 3'h2 == state ? dirty_0_2 : _GEN_8111; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8669 = 3'h2 == state ? dirty_0_3 : _GEN_8112; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8670 = 3'h2 == state ? dirty_0_4 : _GEN_8113; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8671 = 3'h2 == state ? dirty_0_5 : _GEN_8114; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8672 = 3'h2 == state ? dirty_0_6 : _GEN_8115; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8673 = 3'h2 == state ? dirty_0_7 : _GEN_8116; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8674 = 3'h2 == state ? dirty_0_8 : _GEN_8117; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8675 = 3'h2 == state ? dirty_0_9 : _GEN_8118; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8676 = 3'h2 == state ? dirty_0_10 : _GEN_8119; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8677 = 3'h2 == state ? dirty_0_11 : _GEN_8120; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8678 = 3'h2 == state ? dirty_0_12 : _GEN_8121; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8679 = 3'h2 == state ? dirty_0_13 : _GEN_8122; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8680 = 3'h2 == state ? dirty_0_14 : _GEN_8123; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8681 = 3'h2 == state ? dirty_0_15 : _GEN_8124; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8682 = 3'h2 == state ? dirty_0_16 : _GEN_8125; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8683 = 3'h2 == state ? dirty_0_17 : _GEN_8126; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8684 = 3'h2 == state ? dirty_0_18 : _GEN_8127; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8685 = 3'h2 == state ? dirty_0_19 : _GEN_8128; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8686 = 3'h2 == state ? dirty_0_20 : _GEN_8129; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8687 = 3'h2 == state ? dirty_0_21 : _GEN_8130; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8688 = 3'h2 == state ? dirty_0_22 : _GEN_8131; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8689 = 3'h2 == state ? dirty_0_23 : _GEN_8132; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8690 = 3'h2 == state ? dirty_0_24 : _GEN_8133; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8691 = 3'h2 == state ? dirty_0_25 : _GEN_8134; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8692 = 3'h2 == state ? dirty_0_26 : _GEN_8135; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8693 = 3'h2 == state ? dirty_0_27 : _GEN_8136; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8694 = 3'h2 == state ? dirty_0_28 : _GEN_8137; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8695 = 3'h2 == state ? dirty_0_29 : _GEN_8138; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8696 = 3'h2 == state ? dirty_0_30 : _GEN_8139; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8697 = 3'h2 == state ? dirty_0_31 : _GEN_8140; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8698 = 3'h2 == state ? dirty_0_32 : _GEN_8141; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8699 = 3'h2 == state ? dirty_0_33 : _GEN_8142; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8700 = 3'h2 == state ? dirty_0_34 : _GEN_8143; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8701 = 3'h2 == state ? dirty_0_35 : _GEN_8144; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8702 = 3'h2 == state ? dirty_0_36 : _GEN_8145; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8703 = 3'h2 == state ? dirty_0_37 : _GEN_8146; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8704 = 3'h2 == state ? dirty_0_38 : _GEN_8147; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8705 = 3'h2 == state ? dirty_0_39 : _GEN_8148; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8706 = 3'h2 == state ? dirty_0_40 : _GEN_8149; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8707 = 3'h2 == state ? dirty_0_41 : _GEN_8150; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8708 = 3'h2 == state ? dirty_0_42 : _GEN_8151; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8709 = 3'h2 == state ? dirty_0_43 : _GEN_8152; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8710 = 3'h2 == state ? dirty_0_44 : _GEN_8153; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8711 = 3'h2 == state ? dirty_0_45 : _GEN_8154; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8712 = 3'h2 == state ? dirty_0_46 : _GEN_8155; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8713 = 3'h2 == state ? dirty_0_47 : _GEN_8156; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8714 = 3'h2 == state ? dirty_0_48 : _GEN_8157; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8715 = 3'h2 == state ? dirty_0_49 : _GEN_8158; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8716 = 3'h2 == state ? dirty_0_50 : _GEN_8159; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8717 = 3'h2 == state ? dirty_0_51 : _GEN_8160; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8718 = 3'h2 == state ? dirty_0_52 : _GEN_8161; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8719 = 3'h2 == state ? dirty_0_53 : _GEN_8162; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8720 = 3'h2 == state ? dirty_0_54 : _GEN_8163; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8721 = 3'h2 == state ? dirty_0_55 : _GEN_8164; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8722 = 3'h2 == state ? dirty_0_56 : _GEN_8165; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8723 = 3'h2 == state ? dirty_0_57 : _GEN_8166; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8724 = 3'h2 == state ? dirty_0_58 : _GEN_8167; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8725 = 3'h2 == state ? dirty_0_59 : _GEN_8168; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8726 = 3'h2 == state ? dirty_0_60 : _GEN_8169; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8727 = 3'h2 == state ? dirty_0_61 : _GEN_8170; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8728 = 3'h2 == state ? dirty_0_62 : _GEN_8171; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8729 = 3'h2 == state ? dirty_0_63 : _GEN_8172; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8730 = 3'h2 == state ? dirty_0_64 : _GEN_8173; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8731 = 3'h2 == state ? dirty_0_65 : _GEN_8174; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8732 = 3'h2 == state ? dirty_0_66 : _GEN_8175; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8733 = 3'h2 == state ? dirty_0_67 : _GEN_8176; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8734 = 3'h2 == state ? dirty_0_68 : _GEN_8177; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8735 = 3'h2 == state ? dirty_0_69 : _GEN_8178; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8736 = 3'h2 == state ? dirty_0_70 : _GEN_8179; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8737 = 3'h2 == state ? dirty_0_71 : _GEN_8180; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8738 = 3'h2 == state ? dirty_0_72 : _GEN_8181; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8739 = 3'h2 == state ? dirty_0_73 : _GEN_8182; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8740 = 3'h2 == state ? dirty_0_74 : _GEN_8183; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8741 = 3'h2 == state ? dirty_0_75 : _GEN_8184; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8742 = 3'h2 == state ? dirty_0_76 : _GEN_8185; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8743 = 3'h2 == state ? dirty_0_77 : _GEN_8186; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8744 = 3'h2 == state ? dirty_0_78 : _GEN_8187; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8745 = 3'h2 == state ? dirty_0_79 : _GEN_8188; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8746 = 3'h2 == state ? dirty_0_80 : _GEN_8189; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8747 = 3'h2 == state ? dirty_0_81 : _GEN_8190; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8748 = 3'h2 == state ? dirty_0_82 : _GEN_8191; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8749 = 3'h2 == state ? dirty_0_83 : _GEN_8192; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8750 = 3'h2 == state ? dirty_0_84 : _GEN_8193; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8751 = 3'h2 == state ? dirty_0_85 : _GEN_8194; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8752 = 3'h2 == state ? dirty_0_86 : _GEN_8195; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8753 = 3'h2 == state ? dirty_0_87 : _GEN_8196; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8754 = 3'h2 == state ? dirty_0_88 : _GEN_8197; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8755 = 3'h2 == state ? dirty_0_89 : _GEN_8198; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8756 = 3'h2 == state ? dirty_0_90 : _GEN_8199; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8757 = 3'h2 == state ? dirty_0_91 : _GEN_8200; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8758 = 3'h2 == state ? dirty_0_92 : _GEN_8201; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8759 = 3'h2 == state ? dirty_0_93 : _GEN_8202; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8760 = 3'h2 == state ? dirty_0_94 : _GEN_8203; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8761 = 3'h2 == state ? dirty_0_95 : _GEN_8204; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8762 = 3'h2 == state ? dirty_0_96 : _GEN_8205; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8763 = 3'h2 == state ? dirty_0_97 : _GEN_8206; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8764 = 3'h2 == state ? dirty_0_98 : _GEN_8207; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8765 = 3'h2 == state ? dirty_0_99 : _GEN_8208; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8766 = 3'h2 == state ? dirty_0_100 : _GEN_8209; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8767 = 3'h2 == state ? dirty_0_101 : _GEN_8210; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8768 = 3'h2 == state ? dirty_0_102 : _GEN_8211; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8769 = 3'h2 == state ? dirty_0_103 : _GEN_8212; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8770 = 3'h2 == state ? dirty_0_104 : _GEN_8213; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8771 = 3'h2 == state ? dirty_0_105 : _GEN_8214; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8772 = 3'h2 == state ? dirty_0_106 : _GEN_8215; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8773 = 3'h2 == state ? dirty_0_107 : _GEN_8216; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8774 = 3'h2 == state ? dirty_0_108 : _GEN_8217; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8775 = 3'h2 == state ? dirty_0_109 : _GEN_8218; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8776 = 3'h2 == state ? dirty_0_110 : _GEN_8219; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8777 = 3'h2 == state ? dirty_0_111 : _GEN_8220; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8778 = 3'h2 == state ? dirty_0_112 : _GEN_8221; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8779 = 3'h2 == state ? dirty_0_113 : _GEN_8222; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8780 = 3'h2 == state ? dirty_0_114 : _GEN_8223; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8781 = 3'h2 == state ? dirty_0_115 : _GEN_8224; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8782 = 3'h2 == state ? dirty_0_116 : _GEN_8225; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8783 = 3'h2 == state ? dirty_0_117 : _GEN_8226; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8784 = 3'h2 == state ? dirty_0_118 : _GEN_8227; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8785 = 3'h2 == state ? dirty_0_119 : _GEN_8228; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8786 = 3'h2 == state ? dirty_0_120 : _GEN_8229; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8787 = 3'h2 == state ? dirty_0_121 : _GEN_8230; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8788 = 3'h2 == state ? dirty_0_122 : _GEN_8231; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8789 = 3'h2 == state ? dirty_0_123 : _GEN_8232; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8790 = 3'h2 == state ? dirty_0_124 : _GEN_8233; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8791 = 3'h2 == state ? dirty_0_125 : _GEN_8234; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8792 = 3'h2 == state ? dirty_0_126 : _GEN_8235; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8793 = 3'h2 == state ? dirty_0_127 : _GEN_8236; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8794 = 3'h2 == state ? dirty_0_128 : _GEN_8237; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8795 = 3'h2 == state ? dirty_0_129 : _GEN_8238; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8796 = 3'h2 == state ? dirty_0_130 : _GEN_8239; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8797 = 3'h2 == state ? dirty_0_131 : _GEN_8240; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8798 = 3'h2 == state ? dirty_0_132 : _GEN_8241; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8799 = 3'h2 == state ? dirty_0_133 : _GEN_8242; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8800 = 3'h2 == state ? dirty_0_134 : _GEN_8243; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8801 = 3'h2 == state ? dirty_0_135 : _GEN_8244; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8802 = 3'h2 == state ? dirty_0_136 : _GEN_8245; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8803 = 3'h2 == state ? dirty_0_137 : _GEN_8246; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8804 = 3'h2 == state ? dirty_0_138 : _GEN_8247; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8805 = 3'h2 == state ? dirty_0_139 : _GEN_8248; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8806 = 3'h2 == state ? dirty_0_140 : _GEN_8249; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8807 = 3'h2 == state ? dirty_0_141 : _GEN_8250; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8808 = 3'h2 == state ? dirty_0_142 : _GEN_8251; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8809 = 3'h2 == state ? dirty_0_143 : _GEN_8252; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8810 = 3'h2 == state ? dirty_0_144 : _GEN_8253; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8811 = 3'h2 == state ? dirty_0_145 : _GEN_8254; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8812 = 3'h2 == state ? dirty_0_146 : _GEN_8255; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8813 = 3'h2 == state ? dirty_0_147 : _GEN_8256; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8814 = 3'h2 == state ? dirty_0_148 : _GEN_8257; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8815 = 3'h2 == state ? dirty_0_149 : _GEN_8258; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8816 = 3'h2 == state ? dirty_0_150 : _GEN_8259; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8817 = 3'h2 == state ? dirty_0_151 : _GEN_8260; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8818 = 3'h2 == state ? dirty_0_152 : _GEN_8261; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8819 = 3'h2 == state ? dirty_0_153 : _GEN_8262; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8820 = 3'h2 == state ? dirty_0_154 : _GEN_8263; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8821 = 3'h2 == state ? dirty_0_155 : _GEN_8264; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8822 = 3'h2 == state ? dirty_0_156 : _GEN_8265; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8823 = 3'h2 == state ? dirty_0_157 : _GEN_8266; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8824 = 3'h2 == state ? dirty_0_158 : _GEN_8267; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8825 = 3'h2 == state ? dirty_0_159 : _GEN_8268; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8826 = 3'h2 == state ? dirty_0_160 : _GEN_8269; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8827 = 3'h2 == state ? dirty_0_161 : _GEN_8270; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8828 = 3'h2 == state ? dirty_0_162 : _GEN_8271; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8829 = 3'h2 == state ? dirty_0_163 : _GEN_8272; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8830 = 3'h2 == state ? dirty_0_164 : _GEN_8273; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8831 = 3'h2 == state ? dirty_0_165 : _GEN_8274; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8832 = 3'h2 == state ? dirty_0_166 : _GEN_8275; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8833 = 3'h2 == state ? dirty_0_167 : _GEN_8276; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8834 = 3'h2 == state ? dirty_0_168 : _GEN_8277; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8835 = 3'h2 == state ? dirty_0_169 : _GEN_8278; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8836 = 3'h2 == state ? dirty_0_170 : _GEN_8279; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8837 = 3'h2 == state ? dirty_0_171 : _GEN_8280; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8838 = 3'h2 == state ? dirty_0_172 : _GEN_8281; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8839 = 3'h2 == state ? dirty_0_173 : _GEN_8282; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8840 = 3'h2 == state ? dirty_0_174 : _GEN_8283; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8841 = 3'h2 == state ? dirty_0_175 : _GEN_8284; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8842 = 3'h2 == state ? dirty_0_176 : _GEN_8285; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8843 = 3'h2 == state ? dirty_0_177 : _GEN_8286; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8844 = 3'h2 == state ? dirty_0_178 : _GEN_8287; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8845 = 3'h2 == state ? dirty_0_179 : _GEN_8288; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8846 = 3'h2 == state ? dirty_0_180 : _GEN_8289; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8847 = 3'h2 == state ? dirty_0_181 : _GEN_8290; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8848 = 3'h2 == state ? dirty_0_182 : _GEN_8291; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8849 = 3'h2 == state ? dirty_0_183 : _GEN_8292; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8850 = 3'h2 == state ? dirty_0_184 : _GEN_8293; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8851 = 3'h2 == state ? dirty_0_185 : _GEN_8294; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8852 = 3'h2 == state ? dirty_0_186 : _GEN_8295; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8853 = 3'h2 == state ? dirty_0_187 : _GEN_8296; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8854 = 3'h2 == state ? dirty_0_188 : _GEN_8297; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8855 = 3'h2 == state ? dirty_0_189 : _GEN_8298; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8856 = 3'h2 == state ? dirty_0_190 : _GEN_8299; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8857 = 3'h2 == state ? dirty_0_191 : _GEN_8300; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8858 = 3'h2 == state ? dirty_0_192 : _GEN_8301; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8859 = 3'h2 == state ? dirty_0_193 : _GEN_8302; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8860 = 3'h2 == state ? dirty_0_194 : _GEN_8303; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8861 = 3'h2 == state ? dirty_0_195 : _GEN_8304; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8862 = 3'h2 == state ? dirty_0_196 : _GEN_8305; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8863 = 3'h2 == state ? dirty_0_197 : _GEN_8306; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8864 = 3'h2 == state ? dirty_0_198 : _GEN_8307; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8865 = 3'h2 == state ? dirty_0_199 : _GEN_8308; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8866 = 3'h2 == state ? dirty_0_200 : _GEN_8309; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8867 = 3'h2 == state ? dirty_0_201 : _GEN_8310; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8868 = 3'h2 == state ? dirty_0_202 : _GEN_8311; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8869 = 3'h2 == state ? dirty_0_203 : _GEN_8312; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8870 = 3'h2 == state ? dirty_0_204 : _GEN_8313; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8871 = 3'h2 == state ? dirty_0_205 : _GEN_8314; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8872 = 3'h2 == state ? dirty_0_206 : _GEN_8315; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8873 = 3'h2 == state ? dirty_0_207 : _GEN_8316; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8874 = 3'h2 == state ? dirty_0_208 : _GEN_8317; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8875 = 3'h2 == state ? dirty_0_209 : _GEN_8318; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8876 = 3'h2 == state ? dirty_0_210 : _GEN_8319; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8877 = 3'h2 == state ? dirty_0_211 : _GEN_8320; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8878 = 3'h2 == state ? dirty_0_212 : _GEN_8321; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8879 = 3'h2 == state ? dirty_0_213 : _GEN_8322; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8880 = 3'h2 == state ? dirty_0_214 : _GEN_8323; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8881 = 3'h2 == state ? dirty_0_215 : _GEN_8324; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8882 = 3'h2 == state ? dirty_0_216 : _GEN_8325; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8883 = 3'h2 == state ? dirty_0_217 : _GEN_8326; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8884 = 3'h2 == state ? dirty_0_218 : _GEN_8327; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8885 = 3'h2 == state ? dirty_0_219 : _GEN_8328; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8886 = 3'h2 == state ? dirty_0_220 : _GEN_8329; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8887 = 3'h2 == state ? dirty_0_221 : _GEN_8330; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8888 = 3'h2 == state ? dirty_0_222 : _GEN_8331; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8889 = 3'h2 == state ? dirty_0_223 : _GEN_8332; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8890 = 3'h2 == state ? dirty_0_224 : _GEN_8333; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8891 = 3'h2 == state ? dirty_0_225 : _GEN_8334; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8892 = 3'h2 == state ? dirty_0_226 : _GEN_8335; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8893 = 3'h2 == state ? dirty_0_227 : _GEN_8336; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8894 = 3'h2 == state ? dirty_0_228 : _GEN_8337; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8895 = 3'h2 == state ? dirty_0_229 : _GEN_8338; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8896 = 3'h2 == state ? dirty_0_230 : _GEN_8339; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8897 = 3'h2 == state ? dirty_0_231 : _GEN_8340; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8898 = 3'h2 == state ? dirty_0_232 : _GEN_8341; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8899 = 3'h2 == state ? dirty_0_233 : _GEN_8342; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8900 = 3'h2 == state ? dirty_0_234 : _GEN_8343; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8901 = 3'h2 == state ? dirty_0_235 : _GEN_8344; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8902 = 3'h2 == state ? dirty_0_236 : _GEN_8345; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8903 = 3'h2 == state ? dirty_0_237 : _GEN_8346; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8904 = 3'h2 == state ? dirty_0_238 : _GEN_8347; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8905 = 3'h2 == state ? dirty_0_239 : _GEN_8348; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8906 = 3'h2 == state ? dirty_0_240 : _GEN_8349; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8907 = 3'h2 == state ? dirty_0_241 : _GEN_8350; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8908 = 3'h2 == state ? dirty_0_242 : _GEN_8351; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8909 = 3'h2 == state ? dirty_0_243 : _GEN_8352; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8910 = 3'h2 == state ? dirty_0_244 : _GEN_8353; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8911 = 3'h2 == state ? dirty_0_245 : _GEN_8354; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8912 = 3'h2 == state ? dirty_0_246 : _GEN_8355; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8913 = 3'h2 == state ? dirty_0_247 : _GEN_8356; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8914 = 3'h2 == state ? dirty_0_248 : _GEN_8357; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8915 = 3'h2 == state ? dirty_0_249 : _GEN_8358; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8916 = 3'h2 == state ? dirty_0_250 : _GEN_8359; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8917 = 3'h2 == state ? dirty_0_251 : _GEN_8360; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8918 = 3'h2 == state ? dirty_0_252 : _GEN_8361; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8919 = 3'h2 == state ? dirty_0_253 : _GEN_8362; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8920 = 3'h2 == state ? dirty_0_254 : _GEN_8363; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8921 = 3'h2 == state ? dirty_0_255 : _GEN_8364; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8922 = 3'h2 == state ? dirty_1_0 : _GEN_8365; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8923 = 3'h2 == state ? dirty_1_1 : _GEN_8366; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8924 = 3'h2 == state ? dirty_1_2 : _GEN_8367; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8925 = 3'h2 == state ? dirty_1_3 : _GEN_8368; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8926 = 3'h2 == state ? dirty_1_4 : _GEN_8369; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8927 = 3'h2 == state ? dirty_1_5 : _GEN_8370; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8928 = 3'h2 == state ? dirty_1_6 : _GEN_8371; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8929 = 3'h2 == state ? dirty_1_7 : _GEN_8372; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8930 = 3'h2 == state ? dirty_1_8 : _GEN_8373; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8931 = 3'h2 == state ? dirty_1_9 : _GEN_8374; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8932 = 3'h2 == state ? dirty_1_10 : _GEN_8375; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8933 = 3'h2 == state ? dirty_1_11 : _GEN_8376; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8934 = 3'h2 == state ? dirty_1_12 : _GEN_8377; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8935 = 3'h2 == state ? dirty_1_13 : _GEN_8378; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8936 = 3'h2 == state ? dirty_1_14 : _GEN_8379; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8937 = 3'h2 == state ? dirty_1_15 : _GEN_8380; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8938 = 3'h2 == state ? dirty_1_16 : _GEN_8381; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8939 = 3'h2 == state ? dirty_1_17 : _GEN_8382; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8940 = 3'h2 == state ? dirty_1_18 : _GEN_8383; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8941 = 3'h2 == state ? dirty_1_19 : _GEN_8384; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8942 = 3'h2 == state ? dirty_1_20 : _GEN_8385; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8943 = 3'h2 == state ? dirty_1_21 : _GEN_8386; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8944 = 3'h2 == state ? dirty_1_22 : _GEN_8387; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8945 = 3'h2 == state ? dirty_1_23 : _GEN_8388; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8946 = 3'h2 == state ? dirty_1_24 : _GEN_8389; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8947 = 3'h2 == state ? dirty_1_25 : _GEN_8390; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8948 = 3'h2 == state ? dirty_1_26 : _GEN_8391; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8949 = 3'h2 == state ? dirty_1_27 : _GEN_8392; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8950 = 3'h2 == state ? dirty_1_28 : _GEN_8393; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8951 = 3'h2 == state ? dirty_1_29 : _GEN_8394; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8952 = 3'h2 == state ? dirty_1_30 : _GEN_8395; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8953 = 3'h2 == state ? dirty_1_31 : _GEN_8396; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8954 = 3'h2 == state ? dirty_1_32 : _GEN_8397; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8955 = 3'h2 == state ? dirty_1_33 : _GEN_8398; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8956 = 3'h2 == state ? dirty_1_34 : _GEN_8399; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8957 = 3'h2 == state ? dirty_1_35 : _GEN_8400; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8958 = 3'h2 == state ? dirty_1_36 : _GEN_8401; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8959 = 3'h2 == state ? dirty_1_37 : _GEN_8402; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8960 = 3'h2 == state ? dirty_1_38 : _GEN_8403; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8961 = 3'h2 == state ? dirty_1_39 : _GEN_8404; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8962 = 3'h2 == state ? dirty_1_40 : _GEN_8405; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8963 = 3'h2 == state ? dirty_1_41 : _GEN_8406; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8964 = 3'h2 == state ? dirty_1_42 : _GEN_8407; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8965 = 3'h2 == state ? dirty_1_43 : _GEN_8408; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8966 = 3'h2 == state ? dirty_1_44 : _GEN_8409; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8967 = 3'h2 == state ? dirty_1_45 : _GEN_8410; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8968 = 3'h2 == state ? dirty_1_46 : _GEN_8411; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8969 = 3'h2 == state ? dirty_1_47 : _GEN_8412; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8970 = 3'h2 == state ? dirty_1_48 : _GEN_8413; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8971 = 3'h2 == state ? dirty_1_49 : _GEN_8414; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8972 = 3'h2 == state ? dirty_1_50 : _GEN_8415; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8973 = 3'h2 == state ? dirty_1_51 : _GEN_8416; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8974 = 3'h2 == state ? dirty_1_52 : _GEN_8417; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8975 = 3'h2 == state ? dirty_1_53 : _GEN_8418; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8976 = 3'h2 == state ? dirty_1_54 : _GEN_8419; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8977 = 3'h2 == state ? dirty_1_55 : _GEN_8420; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8978 = 3'h2 == state ? dirty_1_56 : _GEN_8421; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8979 = 3'h2 == state ? dirty_1_57 : _GEN_8422; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8980 = 3'h2 == state ? dirty_1_58 : _GEN_8423; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8981 = 3'h2 == state ? dirty_1_59 : _GEN_8424; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8982 = 3'h2 == state ? dirty_1_60 : _GEN_8425; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8983 = 3'h2 == state ? dirty_1_61 : _GEN_8426; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8984 = 3'h2 == state ? dirty_1_62 : _GEN_8427; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8985 = 3'h2 == state ? dirty_1_63 : _GEN_8428; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8986 = 3'h2 == state ? dirty_1_64 : _GEN_8429; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8987 = 3'h2 == state ? dirty_1_65 : _GEN_8430; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8988 = 3'h2 == state ? dirty_1_66 : _GEN_8431; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8989 = 3'h2 == state ? dirty_1_67 : _GEN_8432; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8990 = 3'h2 == state ? dirty_1_68 : _GEN_8433; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8991 = 3'h2 == state ? dirty_1_69 : _GEN_8434; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8992 = 3'h2 == state ? dirty_1_70 : _GEN_8435; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8993 = 3'h2 == state ? dirty_1_71 : _GEN_8436; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8994 = 3'h2 == state ? dirty_1_72 : _GEN_8437; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8995 = 3'h2 == state ? dirty_1_73 : _GEN_8438; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8996 = 3'h2 == state ? dirty_1_74 : _GEN_8439; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8997 = 3'h2 == state ? dirty_1_75 : _GEN_8440; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8998 = 3'h2 == state ? dirty_1_76 : _GEN_8441; // @[dcache.scala 183:18 113:28]
  wire  _GEN_8999 = 3'h2 == state ? dirty_1_77 : _GEN_8442; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9000 = 3'h2 == state ? dirty_1_78 : _GEN_8443; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9001 = 3'h2 == state ? dirty_1_79 : _GEN_8444; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9002 = 3'h2 == state ? dirty_1_80 : _GEN_8445; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9003 = 3'h2 == state ? dirty_1_81 : _GEN_8446; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9004 = 3'h2 == state ? dirty_1_82 : _GEN_8447; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9005 = 3'h2 == state ? dirty_1_83 : _GEN_8448; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9006 = 3'h2 == state ? dirty_1_84 : _GEN_8449; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9007 = 3'h2 == state ? dirty_1_85 : _GEN_8450; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9008 = 3'h2 == state ? dirty_1_86 : _GEN_8451; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9009 = 3'h2 == state ? dirty_1_87 : _GEN_8452; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9010 = 3'h2 == state ? dirty_1_88 : _GEN_8453; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9011 = 3'h2 == state ? dirty_1_89 : _GEN_8454; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9012 = 3'h2 == state ? dirty_1_90 : _GEN_8455; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9013 = 3'h2 == state ? dirty_1_91 : _GEN_8456; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9014 = 3'h2 == state ? dirty_1_92 : _GEN_8457; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9015 = 3'h2 == state ? dirty_1_93 : _GEN_8458; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9016 = 3'h2 == state ? dirty_1_94 : _GEN_8459; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9017 = 3'h2 == state ? dirty_1_95 : _GEN_8460; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9018 = 3'h2 == state ? dirty_1_96 : _GEN_8461; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9019 = 3'h2 == state ? dirty_1_97 : _GEN_8462; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9020 = 3'h2 == state ? dirty_1_98 : _GEN_8463; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9021 = 3'h2 == state ? dirty_1_99 : _GEN_8464; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9022 = 3'h2 == state ? dirty_1_100 : _GEN_8465; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9023 = 3'h2 == state ? dirty_1_101 : _GEN_8466; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9024 = 3'h2 == state ? dirty_1_102 : _GEN_8467; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9025 = 3'h2 == state ? dirty_1_103 : _GEN_8468; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9026 = 3'h2 == state ? dirty_1_104 : _GEN_8469; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9027 = 3'h2 == state ? dirty_1_105 : _GEN_8470; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9028 = 3'h2 == state ? dirty_1_106 : _GEN_8471; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9029 = 3'h2 == state ? dirty_1_107 : _GEN_8472; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9030 = 3'h2 == state ? dirty_1_108 : _GEN_8473; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9031 = 3'h2 == state ? dirty_1_109 : _GEN_8474; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9032 = 3'h2 == state ? dirty_1_110 : _GEN_8475; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9033 = 3'h2 == state ? dirty_1_111 : _GEN_8476; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9034 = 3'h2 == state ? dirty_1_112 : _GEN_8477; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9035 = 3'h2 == state ? dirty_1_113 : _GEN_8478; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9036 = 3'h2 == state ? dirty_1_114 : _GEN_8479; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9037 = 3'h2 == state ? dirty_1_115 : _GEN_8480; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9038 = 3'h2 == state ? dirty_1_116 : _GEN_8481; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9039 = 3'h2 == state ? dirty_1_117 : _GEN_8482; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9040 = 3'h2 == state ? dirty_1_118 : _GEN_8483; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9041 = 3'h2 == state ? dirty_1_119 : _GEN_8484; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9042 = 3'h2 == state ? dirty_1_120 : _GEN_8485; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9043 = 3'h2 == state ? dirty_1_121 : _GEN_8486; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9044 = 3'h2 == state ? dirty_1_122 : _GEN_8487; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9045 = 3'h2 == state ? dirty_1_123 : _GEN_8488; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9046 = 3'h2 == state ? dirty_1_124 : _GEN_8489; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9047 = 3'h2 == state ? dirty_1_125 : _GEN_8490; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9048 = 3'h2 == state ? dirty_1_126 : _GEN_8491; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9049 = 3'h2 == state ? dirty_1_127 : _GEN_8492; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9050 = 3'h2 == state ? dirty_1_128 : _GEN_8493; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9051 = 3'h2 == state ? dirty_1_129 : _GEN_8494; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9052 = 3'h2 == state ? dirty_1_130 : _GEN_8495; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9053 = 3'h2 == state ? dirty_1_131 : _GEN_8496; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9054 = 3'h2 == state ? dirty_1_132 : _GEN_8497; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9055 = 3'h2 == state ? dirty_1_133 : _GEN_8498; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9056 = 3'h2 == state ? dirty_1_134 : _GEN_8499; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9057 = 3'h2 == state ? dirty_1_135 : _GEN_8500; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9058 = 3'h2 == state ? dirty_1_136 : _GEN_8501; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9059 = 3'h2 == state ? dirty_1_137 : _GEN_8502; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9060 = 3'h2 == state ? dirty_1_138 : _GEN_8503; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9061 = 3'h2 == state ? dirty_1_139 : _GEN_8504; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9062 = 3'h2 == state ? dirty_1_140 : _GEN_8505; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9063 = 3'h2 == state ? dirty_1_141 : _GEN_8506; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9064 = 3'h2 == state ? dirty_1_142 : _GEN_8507; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9065 = 3'h2 == state ? dirty_1_143 : _GEN_8508; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9066 = 3'h2 == state ? dirty_1_144 : _GEN_8509; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9067 = 3'h2 == state ? dirty_1_145 : _GEN_8510; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9068 = 3'h2 == state ? dirty_1_146 : _GEN_8511; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9069 = 3'h2 == state ? dirty_1_147 : _GEN_8512; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9070 = 3'h2 == state ? dirty_1_148 : _GEN_8513; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9071 = 3'h2 == state ? dirty_1_149 : _GEN_8514; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9072 = 3'h2 == state ? dirty_1_150 : _GEN_8515; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9073 = 3'h2 == state ? dirty_1_151 : _GEN_8516; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9074 = 3'h2 == state ? dirty_1_152 : _GEN_8517; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9075 = 3'h2 == state ? dirty_1_153 : _GEN_8518; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9076 = 3'h2 == state ? dirty_1_154 : _GEN_8519; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9077 = 3'h2 == state ? dirty_1_155 : _GEN_8520; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9078 = 3'h2 == state ? dirty_1_156 : _GEN_8521; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9079 = 3'h2 == state ? dirty_1_157 : _GEN_8522; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9080 = 3'h2 == state ? dirty_1_158 : _GEN_8523; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9081 = 3'h2 == state ? dirty_1_159 : _GEN_8524; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9082 = 3'h2 == state ? dirty_1_160 : _GEN_8525; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9083 = 3'h2 == state ? dirty_1_161 : _GEN_8526; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9084 = 3'h2 == state ? dirty_1_162 : _GEN_8527; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9085 = 3'h2 == state ? dirty_1_163 : _GEN_8528; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9086 = 3'h2 == state ? dirty_1_164 : _GEN_8529; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9087 = 3'h2 == state ? dirty_1_165 : _GEN_8530; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9088 = 3'h2 == state ? dirty_1_166 : _GEN_8531; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9089 = 3'h2 == state ? dirty_1_167 : _GEN_8532; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9090 = 3'h2 == state ? dirty_1_168 : _GEN_8533; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9091 = 3'h2 == state ? dirty_1_169 : _GEN_8534; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9092 = 3'h2 == state ? dirty_1_170 : _GEN_8535; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9093 = 3'h2 == state ? dirty_1_171 : _GEN_8536; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9094 = 3'h2 == state ? dirty_1_172 : _GEN_8537; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9095 = 3'h2 == state ? dirty_1_173 : _GEN_8538; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9096 = 3'h2 == state ? dirty_1_174 : _GEN_8539; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9097 = 3'h2 == state ? dirty_1_175 : _GEN_8540; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9098 = 3'h2 == state ? dirty_1_176 : _GEN_8541; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9099 = 3'h2 == state ? dirty_1_177 : _GEN_8542; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9100 = 3'h2 == state ? dirty_1_178 : _GEN_8543; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9101 = 3'h2 == state ? dirty_1_179 : _GEN_8544; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9102 = 3'h2 == state ? dirty_1_180 : _GEN_8545; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9103 = 3'h2 == state ? dirty_1_181 : _GEN_8546; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9104 = 3'h2 == state ? dirty_1_182 : _GEN_8547; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9105 = 3'h2 == state ? dirty_1_183 : _GEN_8548; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9106 = 3'h2 == state ? dirty_1_184 : _GEN_8549; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9107 = 3'h2 == state ? dirty_1_185 : _GEN_8550; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9108 = 3'h2 == state ? dirty_1_186 : _GEN_8551; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9109 = 3'h2 == state ? dirty_1_187 : _GEN_8552; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9110 = 3'h2 == state ? dirty_1_188 : _GEN_8553; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9111 = 3'h2 == state ? dirty_1_189 : _GEN_8554; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9112 = 3'h2 == state ? dirty_1_190 : _GEN_8555; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9113 = 3'h2 == state ? dirty_1_191 : _GEN_8556; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9114 = 3'h2 == state ? dirty_1_192 : _GEN_8557; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9115 = 3'h2 == state ? dirty_1_193 : _GEN_8558; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9116 = 3'h2 == state ? dirty_1_194 : _GEN_8559; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9117 = 3'h2 == state ? dirty_1_195 : _GEN_8560; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9118 = 3'h2 == state ? dirty_1_196 : _GEN_8561; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9119 = 3'h2 == state ? dirty_1_197 : _GEN_8562; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9120 = 3'h2 == state ? dirty_1_198 : _GEN_8563; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9121 = 3'h2 == state ? dirty_1_199 : _GEN_8564; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9122 = 3'h2 == state ? dirty_1_200 : _GEN_8565; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9123 = 3'h2 == state ? dirty_1_201 : _GEN_8566; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9124 = 3'h2 == state ? dirty_1_202 : _GEN_8567; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9125 = 3'h2 == state ? dirty_1_203 : _GEN_8568; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9126 = 3'h2 == state ? dirty_1_204 : _GEN_8569; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9127 = 3'h2 == state ? dirty_1_205 : _GEN_8570; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9128 = 3'h2 == state ? dirty_1_206 : _GEN_8571; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9129 = 3'h2 == state ? dirty_1_207 : _GEN_8572; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9130 = 3'h2 == state ? dirty_1_208 : _GEN_8573; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9131 = 3'h2 == state ? dirty_1_209 : _GEN_8574; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9132 = 3'h2 == state ? dirty_1_210 : _GEN_8575; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9133 = 3'h2 == state ? dirty_1_211 : _GEN_8576; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9134 = 3'h2 == state ? dirty_1_212 : _GEN_8577; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9135 = 3'h2 == state ? dirty_1_213 : _GEN_8578; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9136 = 3'h2 == state ? dirty_1_214 : _GEN_8579; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9137 = 3'h2 == state ? dirty_1_215 : _GEN_8580; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9138 = 3'h2 == state ? dirty_1_216 : _GEN_8581; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9139 = 3'h2 == state ? dirty_1_217 : _GEN_8582; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9140 = 3'h2 == state ? dirty_1_218 : _GEN_8583; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9141 = 3'h2 == state ? dirty_1_219 : _GEN_8584; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9142 = 3'h2 == state ? dirty_1_220 : _GEN_8585; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9143 = 3'h2 == state ? dirty_1_221 : _GEN_8586; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9144 = 3'h2 == state ? dirty_1_222 : _GEN_8587; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9145 = 3'h2 == state ? dirty_1_223 : _GEN_8588; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9146 = 3'h2 == state ? dirty_1_224 : _GEN_8589; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9147 = 3'h2 == state ? dirty_1_225 : _GEN_8590; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9148 = 3'h2 == state ? dirty_1_226 : _GEN_8591; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9149 = 3'h2 == state ? dirty_1_227 : _GEN_8592; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9150 = 3'h2 == state ? dirty_1_228 : _GEN_8593; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9151 = 3'h2 == state ? dirty_1_229 : _GEN_8594; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9152 = 3'h2 == state ? dirty_1_230 : _GEN_8595; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9153 = 3'h2 == state ? dirty_1_231 : _GEN_8596; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9154 = 3'h2 == state ? dirty_1_232 : _GEN_8597; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9155 = 3'h2 == state ? dirty_1_233 : _GEN_8598; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9156 = 3'h2 == state ? dirty_1_234 : _GEN_8599; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9157 = 3'h2 == state ? dirty_1_235 : _GEN_8600; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9158 = 3'h2 == state ? dirty_1_236 : _GEN_8601; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9159 = 3'h2 == state ? dirty_1_237 : _GEN_8602; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9160 = 3'h2 == state ? dirty_1_238 : _GEN_8603; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9161 = 3'h2 == state ? dirty_1_239 : _GEN_8604; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9162 = 3'h2 == state ? dirty_1_240 : _GEN_8605; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9163 = 3'h2 == state ? dirty_1_241 : _GEN_8606; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9164 = 3'h2 == state ? dirty_1_242 : _GEN_8607; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9165 = 3'h2 == state ? dirty_1_243 : _GEN_8608; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9166 = 3'h2 == state ? dirty_1_244 : _GEN_8609; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9167 = 3'h2 == state ? dirty_1_245 : _GEN_8610; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9168 = 3'h2 == state ? dirty_1_246 : _GEN_8611; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9169 = 3'h2 == state ? dirty_1_247 : _GEN_8612; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9170 = 3'h2 == state ? dirty_1_248 : _GEN_8613; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9171 = 3'h2 == state ? dirty_1_249 : _GEN_8614; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9172 = 3'h2 == state ? dirty_1_250 : _GEN_8615; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9173 = 3'h2 == state ? dirty_1_251 : _GEN_8616; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9174 = 3'h2 == state ? dirty_1_252 : _GEN_8617; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9175 = 3'h2 == state ? dirty_1_253 : _GEN_8618; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9176 = 3'h2 == state ? dirty_1_254 : _GEN_8619; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9177 = 3'h2 == state ? dirty_1_255 : _GEN_8620; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9178 = 3'h2 == state ? 1'h0 : _GEN_8621; // @[dcache.scala 183:18 144:25]
  wire  _GEN_9179 = 3'h2 == state ? 1'h0 : _GEN_8622; // @[dcache.scala 183:18 144:25]
  wire [20:0] _GEN_9180 = 3'h2 == state ? 21'h0 : _GEN_8623; // @[dcache.scala 183:18 143:25]
  wire [20:0] _GEN_9181 = 3'h2 == state ? 21'h0 : _GEN_8624; // @[dcache.scala 183:18 143:25]
  wire [31:0] _GEN_9182 = 3'h2 == state ? 32'h7777 : _GEN_8625; // @[dcache.scala 183:18 155:25]
  wire  _GEN_9184 = 3'h2 == state ? 1'h0 : _GEN_8627; // @[dcache.scala 183:18 97:21]
  wire [21:0] _GEN_9185 = 3'h2 == state ? 22'h0 : _GEN_8628; // @[dcache.scala 183:18 98:21]
  wire [31:0] _GEN_9193 = 3'h1 == state ? _GEN_73 : _GEN_9182; // @[dcache.scala 183:18]
  wire  _GEN_9201 = 3'h1 == state ? _GEN_81 : _GEN_8645; // @[dcache.scala 183:18]
  wire  _GEN_9205 = 3'h1 == state ? _GEN_125 : _GEN_9184; // @[dcache.scala 183:18]
  wire  _GEN_9212 = 3'h1 == state & _GEN_132; // @[dcache.scala 183:18 156:25]
  wire [7:0] _GEN_9218 = 3'h1 == state ? _GEN_138 : req_set; // @[dcache.scala 183:18 122:34]
  wire  _GEN_9224 = 3'h1 == state ? 1'h0 : _GEN_8640; // @[dcache.scala 183:18 161:25]
  wire [31:0] _GEN_9225 = 3'h1 == state ? 32'h0 : _GEN_8641; // @[dcache.scala 183:18 163:25]
  wire [127:0] _GEN_9226 = 3'h1 == state ? 128'h0 : _GEN_8642; // @[dcache.scala 183:18 165:25]
  wire [2:0] _GEN_9227 = 3'h1 == state ? 3'h0 : _GEN_8643; // @[dcache.scala 183:18 162:25]
  wire [3:0] _GEN_9228 = 3'h1 == state ? 4'h0 : _GEN_8644; // @[dcache.scala 183:18 164:25]
  wire  _GEN_9229 = 3'h1 == state ? 1'h0 : _GEN_8646; // @[dcache.scala 183:18 158:25]
  wire [2:0] _GEN_9230 = 3'h1 == state ? 3'h0 : _GEN_8647; // @[dcache.scala 183:18 159:25]
  wire [31:0] _GEN_9231 = 3'h1 == state ? 32'h0 : _GEN_8648; // @[dcache.scala 183:18 160:25]
  wire [31:0] _GEN_9233 = 3'h1 == state ? 32'h0 : _GEN_8650; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9234 = 3'h1 == state ? 32'h0 : _GEN_8651; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9235 = 3'h1 == state ? 32'h0 : _GEN_8652; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9236 = 3'h1 == state ? 32'h0 : _GEN_8653; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9237 = 3'h1 == state ? 32'h0 : _GEN_8654; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9238 = 3'h1 == state ? 32'h0 : _GEN_8655; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9239 = 3'h1 == state ? 32'h0 : _GEN_8656; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9240 = 3'h1 == state ? 32'h0 : _GEN_8657; // @[dcache.scala 183:18 149:33]
  wire [3:0] _GEN_9241 = 3'h1 == state ? 4'h0 : _GEN_8658; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9242 = 3'h1 == state ? 4'h0 : _GEN_8659; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9243 = 3'h1 == state ? 4'h0 : _GEN_8660; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9244 = 3'h1 == state ? 4'h0 : _GEN_8661; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9245 = 3'h1 == state ? 4'h0 : _GEN_8662; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9246 = 3'h1 == state ? 4'h0 : _GEN_8663; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9247 = 3'h1 == state ? 4'h0 : _GEN_8664; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9248 = 3'h1 == state ? 4'h0 : _GEN_8665; // @[dcache.scala 183:18 150:33]
  wire  _GEN_9249 = 3'h1 == state ? dirty_0_0 : _GEN_8666; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9250 = 3'h1 == state ? dirty_0_1 : _GEN_8667; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9251 = 3'h1 == state ? dirty_0_2 : _GEN_8668; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9252 = 3'h1 == state ? dirty_0_3 : _GEN_8669; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9253 = 3'h1 == state ? dirty_0_4 : _GEN_8670; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9254 = 3'h1 == state ? dirty_0_5 : _GEN_8671; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9255 = 3'h1 == state ? dirty_0_6 : _GEN_8672; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9256 = 3'h1 == state ? dirty_0_7 : _GEN_8673; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9257 = 3'h1 == state ? dirty_0_8 : _GEN_8674; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9258 = 3'h1 == state ? dirty_0_9 : _GEN_8675; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9259 = 3'h1 == state ? dirty_0_10 : _GEN_8676; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9260 = 3'h1 == state ? dirty_0_11 : _GEN_8677; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9261 = 3'h1 == state ? dirty_0_12 : _GEN_8678; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9262 = 3'h1 == state ? dirty_0_13 : _GEN_8679; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9263 = 3'h1 == state ? dirty_0_14 : _GEN_8680; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9264 = 3'h1 == state ? dirty_0_15 : _GEN_8681; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9265 = 3'h1 == state ? dirty_0_16 : _GEN_8682; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9266 = 3'h1 == state ? dirty_0_17 : _GEN_8683; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9267 = 3'h1 == state ? dirty_0_18 : _GEN_8684; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9268 = 3'h1 == state ? dirty_0_19 : _GEN_8685; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9269 = 3'h1 == state ? dirty_0_20 : _GEN_8686; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9270 = 3'h1 == state ? dirty_0_21 : _GEN_8687; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9271 = 3'h1 == state ? dirty_0_22 : _GEN_8688; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9272 = 3'h1 == state ? dirty_0_23 : _GEN_8689; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9273 = 3'h1 == state ? dirty_0_24 : _GEN_8690; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9274 = 3'h1 == state ? dirty_0_25 : _GEN_8691; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9275 = 3'h1 == state ? dirty_0_26 : _GEN_8692; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9276 = 3'h1 == state ? dirty_0_27 : _GEN_8693; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9277 = 3'h1 == state ? dirty_0_28 : _GEN_8694; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9278 = 3'h1 == state ? dirty_0_29 : _GEN_8695; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9279 = 3'h1 == state ? dirty_0_30 : _GEN_8696; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9280 = 3'h1 == state ? dirty_0_31 : _GEN_8697; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9281 = 3'h1 == state ? dirty_0_32 : _GEN_8698; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9282 = 3'h1 == state ? dirty_0_33 : _GEN_8699; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9283 = 3'h1 == state ? dirty_0_34 : _GEN_8700; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9284 = 3'h1 == state ? dirty_0_35 : _GEN_8701; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9285 = 3'h1 == state ? dirty_0_36 : _GEN_8702; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9286 = 3'h1 == state ? dirty_0_37 : _GEN_8703; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9287 = 3'h1 == state ? dirty_0_38 : _GEN_8704; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9288 = 3'h1 == state ? dirty_0_39 : _GEN_8705; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9289 = 3'h1 == state ? dirty_0_40 : _GEN_8706; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9290 = 3'h1 == state ? dirty_0_41 : _GEN_8707; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9291 = 3'h1 == state ? dirty_0_42 : _GEN_8708; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9292 = 3'h1 == state ? dirty_0_43 : _GEN_8709; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9293 = 3'h1 == state ? dirty_0_44 : _GEN_8710; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9294 = 3'h1 == state ? dirty_0_45 : _GEN_8711; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9295 = 3'h1 == state ? dirty_0_46 : _GEN_8712; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9296 = 3'h1 == state ? dirty_0_47 : _GEN_8713; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9297 = 3'h1 == state ? dirty_0_48 : _GEN_8714; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9298 = 3'h1 == state ? dirty_0_49 : _GEN_8715; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9299 = 3'h1 == state ? dirty_0_50 : _GEN_8716; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9300 = 3'h1 == state ? dirty_0_51 : _GEN_8717; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9301 = 3'h1 == state ? dirty_0_52 : _GEN_8718; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9302 = 3'h1 == state ? dirty_0_53 : _GEN_8719; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9303 = 3'h1 == state ? dirty_0_54 : _GEN_8720; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9304 = 3'h1 == state ? dirty_0_55 : _GEN_8721; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9305 = 3'h1 == state ? dirty_0_56 : _GEN_8722; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9306 = 3'h1 == state ? dirty_0_57 : _GEN_8723; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9307 = 3'h1 == state ? dirty_0_58 : _GEN_8724; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9308 = 3'h1 == state ? dirty_0_59 : _GEN_8725; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9309 = 3'h1 == state ? dirty_0_60 : _GEN_8726; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9310 = 3'h1 == state ? dirty_0_61 : _GEN_8727; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9311 = 3'h1 == state ? dirty_0_62 : _GEN_8728; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9312 = 3'h1 == state ? dirty_0_63 : _GEN_8729; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9313 = 3'h1 == state ? dirty_0_64 : _GEN_8730; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9314 = 3'h1 == state ? dirty_0_65 : _GEN_8731; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9315 = 3'h1 == state ? dirty_0_66 : _GEN_8732; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9316 = 3'h1 == state ? dirty_0_67 : _GEN_8733; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9317 = 3'h1 == state ? dirty_0_68 : _GEN_8734; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9318 = 3'h1 == state ? dirty_0_69 : _GEN_8735; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9319 = 3'h1 == state ? dirty_0_70 : _GEN_8736; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9320 = 3'h1 == state ? dirty_0_71 : _GEN_8737; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9321 = 3'h1 == state ? dirty_0_72 : _GEN_8738; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9322 = 3'h1 == state ? dirty_0_73 : _GEN_8739; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9323 = 3'h1 == state ? dirty_0_74 : _GEN_8740; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9324 = 3'h1 == state ? dirty_0_75 : _GEN_8741; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9325 = 3'h1 == state ? dirty_0_76 : _GEN_8742; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9326 = 3'h1 == state ? dirty_0_77 : _GEN_8743; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9327 = 3'h1 == state ? dirty_0_78 : _GEN_8744; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9328 = 3'h1 == state ? dirty_0_79 : _GEN_8745; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9329 = 3'h1 == state ? dirty_0_80 : _GEN_8746; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9330 = 3'h1 == state ? dirty_0_81 : _GEN_8747; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9331 = 3'h1 == state ? dirty_0_82 : _GEN_8748; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9332 = 3'h1 == state ? dirty_0_83 : _GEN_8749; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9333 = 3'h1 == state ? dirty_0_84 : _GEN_8750; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9334 = 3'h1 == state ? dirty_0_85 : _GEN_8751; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9335 = 3'h1 == state ? dirty_0_86 : _GEN_8752; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9336 = 3'h1 == state ? dirty_0_87 : _GEN_8753; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9337 = 3'h1 == state ? dirty_0_88 : _GEN_8754; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9338 = 3'h1 == state ? dirty_0_89 : _GEN_8755; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9339 = 3'h1 == state ? dirty_0_90 : _GEN_8756; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9340 = 3'h1 == state ? dirty_0_91 : _GEN_8757; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9341 = 3'h1 == state ? dirty_0_92 : _GEN_8758; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9342 = 3'h1 == state ? dirty_0_93 : _GEN_8759; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9343 = 3'h1 == state ? dirty_0_94 : _GEN_8760; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9344 = 3'h1 == state ? dirty_0_95 : _GEN_8761; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9345 = 3'h1 == state ? dirty_0_96 : _GEN_8762; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9346 = 3'h1 == state ? dirty_0_97 : _GEN_8763; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9347 = 3'h1 == state ? dirty_0_98 : _GEN_8764; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9348 = 3'h1 == state ? dirty_0_99 : _GEN_8765; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9349 = 3'h1 == state ? dirty_0_100 : _GEN_8766; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9350 = 3'h1 == state ? dirty_0_101 : _GEN_8767; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9351 = 3'h1 == state ? dirty_0_102 : _GEN_8768; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9352 = 3'h1 == state ? dirty_0_103 : _GEN_8769; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9353 = 3'h1 == state ? dirty_0_104 : _GEN_8770; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9354 = 3'h1 == state ? dirty_0_105 : _GEN_8771; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9355 = 3'h1 == state ? dirty_0_106 : _GEN_8772; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9356 = 3'h1 == state ? dirty_0_107 : _GEN_8773; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9357 = 3'h1 == state ? dirty_0_108 : _GEN_8774; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9358 = 3'h1 == state ? dirty_0_109 : _GEN_8775; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9359 = 3'h1 == state ? dirty_0_110 : _GEN_8776; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9360 = 3'h1 == state ? dirty_0_111 : _GEN_8777; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9361 = 3'h1 == state ? dirty_0_112 : _GEN_8778; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9362 = 3'h1 == state ? dirty_0_113 : _GEN_8779; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9363 = 3'h1 == state ? dirty_0_114 : _GEN_8780; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9364 = 3'h1 == state ? dirty_0_115 : _GEN_8781; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9365 = 3'h1 == state ? dirty_0_116 : _GEN_8782; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9366 = 3'h1 == state ? dirty_0_117 : _GEN_8783; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9367 = 3'h1 == state ? dirty_0_118 : _GEN_8784; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9368 = 3'h1 == state ? dirty_0_119 : _GEN_8785; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9369 = 3'h1 == state ? dirty_0_120 : _GEN_8786; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9370 = 3'h1 == state ? dirty_0_121 : _GEN_8787; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9371 = 3'h1 == state ? dirty_0_122 : _GEN_8788; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9372 = 3'h1 == state ? dirty_0_123 : _GEN_8789; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9373 = 3'h1 == state ? dirty_0_124 : _GEN_8790; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9374 = 3'h1 == state ? dirty_0_125 : _GEN_8791; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9375 = 3'h1 == state ? dirty_0_126 : _GEN_8792; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9376 = 3'h1 == state ? dirty_0_127 : _GEN_8793; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9377 = 3'h1 == state ? dirty_0_128 : _GEN_8794; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9378 = 3'h1 == state ? dirty_0_129 : _GEN_8795; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9379 = 3'h1 == state ? dirty_0_130 : _GEN_8796; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9380 = 3'h1 == state ? dirty_0_131 : _GEN_8797; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9381 = 3'h1 == state ? dirty_0_132 : _GEN_8798; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9382 = 3'h1 == state ? dirty_0_133 : _GEN_8799; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9383 = 3'h1 == state ? dirty_0_134 : _GEN_8800; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9384 = 3'h1 == state ? dirty_0_135 : _GEN_8801; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9385 = 3'h1 == state ? dirty_0_136 : _GEN_8802; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9386 = 3'h1 == state ? dirty_0_137 : _GEN_8803; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9387 = 3'h1 == state ? dirty_0_138 : _GEN_8804; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9388 = 3'h1 == state ? dirty_0_139 : _GEN_8805; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9389 = 3'h1 == state ? dirty_0_140 : _GEN_8806; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9390 = 3'h1 == state ? dirty_0_141 : _GEN_8807; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9391 = 3'h1 == state ? dirty_0_142 : _GEN_8808; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9392 = 3'h1 == state ? dirty_0_143 : _GEN_8809; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9393 = 3'h1 == state ? dirty_0_144 : _GEN_8810; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9394 = 3'h1 == state ? dirty_0_145 : _GEN_8811; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9395 = 3'h1 == state ? dirty_0_146 : _GEN_8812; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9396 = 3'h1 == state ? dirty_0_147 : _GEN_8813; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9397 = 3'h1 == state ? dirty_0_148 : _GEN_8814; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9398 = 3'h1 == state ? dirty_0_149 : _GEN_8815; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9399 = 3'h1 == state ? dirty_0_150 : _GEN_8816; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9400 = 3'h1 == state ? dirty_0_151 : _GEN_8817; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9401 = 3'h1 == state ? dirty_0_152 : _GEN_8818; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9402 = 3'h1 == state ? dirty_0_153 : _GEN_8819; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9403 = 3'h1 == state ? dirty_0_154 : _GEN_8820; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9404 = 3'h1 == state ? dirty_0_155 : _GEN_8821; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9405 = 3'h1 == state ? dirty_0_156 : _GEN_8822; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9406 = 3'h1 == state ? dirty_0_157 : _GEN_8823; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9407 = 3'h1 == state ? dirty_0_158 : _GEN_8824; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9408 = 3'h1 == state ? dirty_0_159 : _GEN_8825; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9409 = 3'h1 == state ? dirty_0_160 : _GEN_8826; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9410 = 3'h1 == state ? dirty_0_161 : _GEN_8827; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9411 = 3'h1 == state ? dirty_0_162 : _GEN_8828; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9412 = 3'h1 == state ? dirty_0_163 : _GEN_8829; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9413 = 3'h1 == state ? dirty_0_164 : _GEN_8830; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9414 = 3'h1 == state ? dirty_0_165 : _GEN_8831; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9415 = 3'h1 == state ? dirty_0_166 : _GEN_8832; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9416 = 3'h1 == state ? dirty_0_167 : _GEN_8833; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9417 = 3'h1 == state ? dirty_0_168 : _GEN_8834; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9418 = 3'h1 == state ? dirty_0_169 : _GEN_8835; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9419 = 3'h1 == state ? dirty_0_170 : _GEN_8836; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9420 = 3'h1 == state ? dirty_0_171 : _GEN_8837; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9421 = 3'h1 == state ? dirty_0_172 : _GEN_8838; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9422 = 3'h1 == state ? dirty_0_173 : _GEN_8839; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9423 = 3'h1 == state ? dirty_0_174 : _GEN_8840; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9424 = 3'h1 == state ? dirty_0_175 : _GEN_8841; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9425 = 3'h1 == state ? dirty_0_176 : _GEN_8842; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9426 = 3'h1 == state ? dirty_0_177 : _GEN_8843; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9427 = 3'h1 == state ? dirty_0_178 : _GEN_8844; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9428 = 3'h1 == state ? dirty_0_179 : _GEN_8845; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9429 = 3'h1 == state ? dirty_0_180 : _GEN_8846; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9430 = 3'h1 == state ? dirty_0_181 : _GEN_8847; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9431 = 3'h1 == state ? dirty_0_182 : _GEN_8848; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9432 = 3'h1 == state ? dirty_0_183 : _GEN_8849; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9433 = 3'h1 == state ? dirty_0_184 : _GEN_8850; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9434 = 3'h1 == state ? dirty_0_185 : _GEN_8851; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9435 = 3'h1 == state ? dirty_0_186 : _GEN_8852; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9436 = 3'h1 == state ? dirty_0_187 : _GEN_8853; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9437 = 3'h1 == state ? dirty_0_188 : _GEN_8854; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9438 = 3'h1 == state ? dirty_0_189 : _GEN_8855; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9439 = 3'h1 == state ? dirty_0_190 : _GEN_8856; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9440 = 3'h1 == state ? dirty_0_191 : _GEN_8857; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9441 = 3'h1 == state ? dirty_0_192 : _GEN_8858; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9442 = 3'h1 == state ? dirty_0_193 : _GEN_8859; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9443 = 3'h1 == state ? dirty_0_194 : _GEN_8860; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9444 = 3'h1 == state ? dirty_0_195 : _GEN_8861; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9445 = 3'h1 == state ? dirty_0_196 : _GEN_8862; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9446 = 3'h1 == state ? dirty_0_197 : _GEN_8863; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9447 = 3'h1 == state ? dirty_0_198 : _GEN_8864; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9448 = 3'h1 == state ? dirty_0_199 : _GEN_8865; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9449 = 3'h1 == state ? dirty_0_200 : _GEN_8866; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9450 = 3'h1 == state ? dirty_0_201 : _GEN_8867; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9451 = 3'h1 == state ? dirty_0_202 : _GEN_8868; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9452 = 3'h1 == state ? dirty_0_203 : _GEN_8869; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9453 = 3'h1 == state ? dirty_0_204 : _GEN_8870; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9454 = 3'h1 == state ? dirty_0_205 : _GEN_8871; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9455 = 3'h1 == state ? dirty_0_206 : _GEN_8872; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9456 = 3'h1 == state ? dirty_0_207 : _GEN_8873; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9457 = 3'h1 == state ? dirty_0_208 : _GEN_8874; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9458 = 3'h1 == state ? dirty_0_209 : _GEN_8875; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9459 = 3'h1 == state ? dirty_0_210 : _GEN_8876; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9460 = 3'h1 == state ? dirty_0_211 : _GEN_8877; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9461 = 3'h1 == state ? dirty_0_212 : _GEN_8878; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9462 = 3'h1 == state ? dirty_0_213 : _GEN_8879; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9463 = 3'h1 == state ? dirty_0_214 : _GEN_8880; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9464 = 3'h1 == state ? dirty_0_215 : _GEN_8881; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9465 = 3'h1 == state ? dirty_0_216 : _GEN_8882; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9466 = 3'h1 == state ? dirty_0_217 : _GEN_8883; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9467 = 3'h1 == state ? dirty_0_218 : _GEN_8884; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9468 = 3'h1 == state ? dirty_0_219 : _GEN_8885; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9469 = 3'h1 == state ? dirty_0_220 : _GEN_8886; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9470 = 3'h1 == state ? dirty_0_221 : _GEN_8887; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9471 = 3'h1 == state ? dirty_0_222 : _GEN_8888; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9472 = 3'h1 == state ? dirty_0_223 : _GEN_8889; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9473 = 3'h1 == state ? dirty_0_224 : _GEN_8890; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9474 = 3'h1 == state ? dirty_0_225 : _GEN_8891; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9475 = 3'h1 == state ? dirty_0_226 : _GEN_8892; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9476 = 3'h1 == state ? dirty_0_227 : _GEN_8893; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9477 = 3'h1 == state ? dirty_0_228 : _GEN_8894; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9478 = 3'h1 == state ? dirty_0_229 : _GEN_8895; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9479 = 3'h1 == state ? dirty_0_230 : _GEN_8896; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9480 = 3'h1 == state ? dirty_0_231 : _GEN_8897; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9481 = 3'h1 == state ? dirty_0_232 : _GEN_8898; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9482 = 3'h1 == state ? dirty_0_233 : _GEN_8899; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9483 = 3'h1 == state ? dirty_0_234 : _GEN_8900; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9484 = 3'h1 == state ? dirty_0_235 : _GEN_8901; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9485 = 3'h1 == state ? dirty_0_236 : _GEN_8902; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9486 = 3'h1 == state ? dirty_0_237 : _GEN_8903; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9487 = 3'h1 == state ? dirty_0_238 : _GEN_8904; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9488 = 3'h1 == state ? dirty_0_239 : _GEN_8905; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9489 = 3'h1 == state ? dirty_0_240 : _GEN_8906; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9490 = 3'h1 == state ? dirty_0_241 : _GEN_8907; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9491 = 3'h1 == state ? dirty_0_242 : _GEN_8908; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9492 = 3'h1 == state ? dirty_0_243 : _GEN_8909; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9493 = 3'h1 == state ? dirty_0_244 : _GEN_8910; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9494 = 3'h1 == state ? dirty_0_245 : _GEN_8911; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9495 = 3'h1 == state ? dirty_0_246 : _GEN_8912; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9496 = 3'h1 == state ? dirty_0_247 : _GEN_8913; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9497 = 3'h1 == state ? dirty_0_248 : _GEN_8914; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9498 = 3'h1 == state ? dirty_0_249 : _GEN_8915; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9499 = 3'h1 == state ? dirty_0_250 : _GEN_8916; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9500 = 3'h1 == state ? dirty_0_251 : _GEN_8917; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9501 = 3'h1 == state ? dirty_0_252 : _GEN_8918; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9502 = 3'h1 == state ? dirty_0_253 : _GEN_8919; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9503 = 3'h1 == state ? dirty_0_254 : _GEN_8920; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9504 = 3'h1 == state ? dirty_0_255 : _GEN_8921; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9505 = 3'h1 == state ? dirty_1_0 : _GEN_8922; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9506 = 3'h1 == state ? dirty_1_1 : _GEN_8923; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9507 = 3'h1 == state ? dirty_1_2 : _GEN_8924; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9508 = 3'h1 == state ? dirty_1_3 : _GEN_8925; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9509 = 3'h1 == state ? dirty_1_4 : _GEN_8926; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9510 = 3'h1 == state ? dirty_1_5 : _GEN_8927; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9511 = 3'h1 == state ? dirty_1_6 : _GEN_8928; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9512 = 3'h1 == state ? dirty_1_7 : _GEN_8929; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9513 = 3'h1 == state ? dirty_1_8 : _GEN_8930; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9514 = 3'h1 == state ? dirty_1_9 : _GEN_8931; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9515 = 3'h1 == state ? dirty_1_10 : _GEN_8932; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9516 = 3'h1 == state ? dirty_1_11 : _GEN_8933; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9517 = 3'h1 == state ? dirty_1_12 : _GEN_8934; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9518 = 3'h1 == state ? dirty_1_13 : _GEN_8935; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9519 = 3'h1 == state ? dirty_1_14 : _GEN_8936; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9520 = 3'h1 == state ? dirty_1_15 : _GEN_8937; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9521 = 3'h1 == state ? dirty_1_16 : _GEN_8938; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9522 = 3'h1 == state ? dirty_1_17 : _GEN_8939; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9523 = 3'h1 == state ? dirty_1_18 : _GEN_8940; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9524 = 3'h1 == state ? dirty_1_19 : _GEN_8941; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9525 = 3'h1 == state ? dirty_1_20 : _GEN_8942; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9526 = 3'h1 == state ? dirty_1_21 : _GEN_8943; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9527 = 3'h1 == state ? dirty_1_22 : _GEN_8944; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9528 = 3'h1 == state ? dirty_1_23 : _GEN_8945; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9529 = 3'h1 == state ? dirty_1_24 : _GEN_8946; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9530 = 3'h1 == state ? dirty_1_25 : _GEN_8947; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9531 = 3'h1 == state ? dirty_1_26 : _GEN_8948; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9532 = 3'h1 == state ? dirty_1_27 : _GEN_8949; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9533 = 3'h1 == state ? dirty_1_28 : _GEN_8950; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9534 = 3'h1 == state ? dirty_1_29 : _GEN_8951; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9535 = 3'h1 == state ? dirty_1_30 : _GEN_8952; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9536 = 3'h1 == state ? dirty_1_31 : _GEN_8953; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9537 = 3'h1 == state ? dirty_1_32 : _GEN_8954; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9538 = 3'h1 == state ? dirty_1_33 : _GEN_8955; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9539 = 3'h1 == state ? dirty_1_34 : _GEN_8956; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9540 = 3'h1 == state ? dirty_1_35 : _GEN_8957; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9541 = 3'h1 == state ? dirty_1_36 : _GEN_8958; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9542 = 3'h1 == state ? dirty_1_37 : _GEN_8959; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9543 = 3'h1 == state ? dirty_1_38 : _GEN_8960; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9544 = 3'h1 == state ? dirty_1_39 : _GEN_8961; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9545 = 3'h1 == state ? dirty_1_40 : _GEN_8962; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9546 = 3'h1 == state ? dirty_1_41 : _GEN_8963; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9547 = 3'h1 == state ? dirty_1_42 : _GEN_8964; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9548 = 3'h1 == state ? dirty_1_43 : _GEN_8965; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9549 = 3'h1 == state ? dirty_1_44 : _GEN_8966; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9550 = 3'h1 == state ? dirty_1_45 : _GEN_8967; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9551 = 3'h1 == state ? dirty_1_46 : _GEN_8968; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9552 = 3'h1 == state ? dirty_1_47 : _GEN_8969; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9553 = 3'h1 == state ? dirty_1_48 : _GEN_8970; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9554 = 3'h1 == state ? dirty_1_49 : _GEN_8971; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9555 = 3'h1 == state ? dirty_1_50 : _GEN_8972; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9556 = 3'h1 == state ? dirty_1_51 : _GEN_8973; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9557 = 3'h1 == state ? dirty_1_52 : _GEN_8974; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9558 = 3'h1 == state ? dirty_1_53 : _GEN_8975; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9559 = 3'h1 == state ? dirty_1_54 : _GEN_8976; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9560 = 3'h1 == state ? dirty_1_55 : _GEN_8977; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9561 = 3'h1 == state ? dirty_1_56 : _GEN_8978; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9562 = 3'h1 == state ? dirty_1_57 : _GEN_8979; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9563 = 3'h1 == state ? dirty_1_58 : _GEN_8980; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9564 = 3'h1 == state ? dirty_1_59 : _GEN_8981; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9565 = 3'h1 == state ? dirty_1_60 : _GEN_8982; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9566 = 3'h1 == state ? dirty_1_61 : _GEN_8983; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9567 = 3'h1 == state ? dirty_1_62 : _GEN_8984; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9568 = 3'h1 == state ? dirty_1_63 : _GEN_8985; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9569 = 3'h1 == state ? dirty_1_64 : _GEN_8986; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9570 = 3'h1 == state ? dirty_1_65 : _GEN_8987; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9571 = 3'h1 == state ? dirty_1_66 : _GEN_8988; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9572 = 3'h1 == state ? dirty_1_67 : _GEN_8989; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9573 = 3'h1 == state ? dirty_1_68 : _GEN_8990; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9574 = 3'h1 == state ? dirty_1_69 : _GEN_8991; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9575 = 3'h1 == state ? dirty_1_70 : _GEN_8992; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9576 = 3'h1 == state ? dirty_1_71 : _GEN_8993; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9577 = 3'h1 == state ? dirty_1_72 : _GEN_8994; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9578 = 3'h1 == state ? dirty_1_73 : _GEN_8995; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9579 = 3'h1 == state ? dirty_1_74 : _GEN_8996; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9580 = 3'h1 == state ? dirty_1_75 : _GEN_8997; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9581 = 3'h1 == state ? dirty_1_76 : _GEN_8998; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9582 = 3'h1 == state ? dirty_1_77 : _GEN_8999; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9583 = 3'h1 == state ? dirty_1_78 : _GEN_9000; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9584 = 3'h1 == state ? dirty_1_79 : _GEN_9001; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9585 = 3'h1 == state ? dirty_1_80 : _GEN_9002; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9586 = 3'h1 == state ? dirty_1_81 : _GEN_9003; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9587 = 3'h1 == state ? dirty_1_82 : _GEN_9004; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9588 = 3'h1 == state ? dirty_1_83 : _GEN_9005; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9589 = 3'h1 == state ? dirty_1_84 : _GEN_9006; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9590 = 3'h1 == state ? dirty_1_85 : _GEN_9007; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9591 = 3'h1 == state ? dirty_1_86 : _GEN_9008; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9592 = 3'h1 == state ? dirty_1_87 : _GEN_9009; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9593 = 3'h1 == state ? dirty_1_88 : _GEN_9010; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9594 = 3'h1 == state ? dirty_1_89 : _GEN_9011; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9595 = 3'h1 == state ? dirty_1_90 : _GEN_9012; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9596 = 3'h1 == state ? dirty_1_91 : _GEN_9013; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9597 = 3'h1 == state ? dirty_1_92 : _GEN_9014; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9598 = 3'h1 == state ? dirty_1_93 : _GEN_9015; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9599 = 3'h1 == state ? dirty_1_94 : _GEN_9016; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9600 = 3'h1 == state ? dirty_1_95 : _GEN_9017; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9601 = 3'h1 == state ? dirty_1_96 : _GEN_9018; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9602 = 3'h1 == state ? dirty_1_97 : _GEN_9019; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9603 = 3'h1 == state ? dirty_1_98 : _GEN_9020; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9604 = 3'h1 == state ? dirty_1_99 : _GEN_9021; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9605 = 3'h1 == state ? dirty_1_100 : _GEN_9022; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9606 = 3'h1 == state ? dirty_1_101 : _GEN_9023; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9607 = 3'h1 == state ? dirty_1_102 : _GEN_9024; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9608 = 3'h1 == state ? dirty_1_103 : _GEN_9025; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9609 = 3'h1 == state ? dirty_1_104 : _GEN_9026; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9610 = 3'h1 == state ? dirty_1_105 : _GEN_9027; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9611 = 3'h1 == state ? dirty_1_106 : _GEN_9028; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9612 = 3'h1 == state ? dirty_1_107 : _GEN_9029; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9613 = 3'h1 == state ? dirty_1_108 : _GEN_9030; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9614 = 3'h1 == state ? dirty_1_109 : _GEN_9031; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9615 = 3'h1 == state ? dirty_1_110 : _GEN_9032; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9616 = 3'h1 == state ? dirty_1_111 : _GEN_9033; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9617 = 3'h1 == state ? dirty_1_112 : _GEN_9034; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9618 = 3'h1 == state ? dirty_1_113 : _GEN_9035; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9619 = 3'h1 == state ? dirty_1_114 : _GEN_9036; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9620 = 3'h1 == state ? dirty_1_115 : _GEN_9037; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9621 = 3'h1 == state ? dirty_1_116 : _GEN_9038; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9622 = 3'h1 == state ? dirty_1_117 : _GEN_9039; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9623 = 3'h1 == state ? dirty_1_118 : _GEN_9040; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9624 = 3'h1 == state ? dirty_1_119 : _GEN_9041; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9625 = 3'h1 == state ? dirty_1_120 : _GEN_9042; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9626 = 3'h1 == state ? dirty_1_121 : _GEN_9043; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9627 = 3'h1 == state ? dirty_1_122 : _GEN_9044; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9628 = 3'h1 == state ? dirty_1_123 : _GEN_9045; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9629 = 3'h1 == state ? dirty_1_124 : _GEN_9046; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9630 = 3'h1 == state ? dirty_1_125 : _GEN_9047; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9631 = 3'h1 == state ? dirty_1_126 : _GEN_9048; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9632 = 3'h1 == state ? dirty_1_127 : _GEN_9049; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9633 = 3'h1 == state ? dirty_1_128 : _GEN_9050; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9634 = 3'h1 == state ? dirty_1_129 : _GEN_9051; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9635 = 3'h1 == state ? dirty_1_130 : _GEN_9052; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9636 = 3'h1 == state ? dirty_1_131 : _GEN_9053; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9637 = 3'h1 == state ? dirty_1_132 : _GEN_9054; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9638 = 3'h1 == state ? dirty_1_133 : _GEN_9055; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9639 = 3'h1 == state ? dirty_1_134 : _GEN_9056; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9640 = 3'h1 == state ? dirty_1_135 : _GEN_9057; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9641 = 3'h1 == state ? dirty_1_136 : _GEN_9058; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9642 = 3'h1 == state ? dirty_1_137 : _GEN_9059; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9643 = 3'h1 == state ? dirty_1_138 : _GEN_9060; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9644 = 3'h1 == state ? dirty_1_139 : _GEN_9061; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9645 = 3'h1 == state ? dirty_1_140 : _GEN_9062; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9646 = 3'h1 == state ? dirty_1_141 : _GEN_9063; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9647 = 3'h1 == state ? dirty_1_142 : _GEN_9064; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9648 = 3'h1 == state ? dirty_1_143 : _GEN_9065; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9649 = 3'h1 == state ? dirty_1_144 : _GEN_9066; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9650 = 3'h1 == state ? dirty_1_145 : _GEN_9067; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9651 = 3'h1 == state ? dirty_1_146 : _GEN_9068; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9652 = 3'h1 == state ? dirty_1_147 : _GEN_9069; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9653 = 3'h1 == state ? dirty_1_148 : _GEN_9070; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9654 = 3'h1 == state ? dirty_1_149 : _GEN_9071; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9655 = 3'h1 == state ? dirty_1_150 : _GEN_9072; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9656 = 3'h1 == state ? dirty_1_151 : _GEN_9073; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9657 = 3'h1 == state ? dirty_1_152 : _GEN_9074; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9658 = 3'h1 == state ? dirty_1_153 : _GEN_9075; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9659 = 3'h1 == state ? dirty_1_154 : _GEN_9076; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9660 = 3'h1 == state ? dirty_1_155 : _GEN_9077; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9661 = 3'h1 == state ? dirty_1_156 : _GEN_9078; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9662 = 3'h1 == state ? dirty_1_157 : _GEN_9079; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9663 = 3'h1 == state ? dirty_1_158 : _GEN_9080; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9664 = 3'h1 == state ? dirty_1_159 : _GEN_9081; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9665 = 3'h1 == state ? dirty_1_160 : _GEN_9082; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9666 = 3'h1 == state ? dirty_1_161 : _GEN_9083; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9667 = 3'h1 == state ? dirty_1_162 : _GEN_9084; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9668 = 3'h1 == state ? dirty_1_163 : _GEN_9085; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9669 = 3'h1 == state ? dirty_1_164 : _GEN_9086; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9670 = 3'h1 == state ? dirty_1_165 : _GEN_9087; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9671 = 3'h1 == state ? dirty_1_166 : _GEN_9088; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9672 = 3'h1 == state ? dirty_1_167 : _GEN_9089; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9673 = 3'h1 == state ? dirty_1_168 : _GEN_9090; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9674 = 3'h1 == state ? dirty_1_169 : _GEN_9091; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9675 = 3'h1 == state ? dirty_1_170 : _GEN_9092; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9676 = 3'h1 == state ? dirty_1_171 : _GEN_9093; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9677 = 3'h1 == state ? dirty_1_172 : _GEN_9094; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9678 = 3'h1 == state ? dirty_1_173 : _GEN_9095; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9679 = 3'h1 == state ? dirty_1_174 : _GEN_9096; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9680 = 3'h1 == state ? dirty_1_175 : _GEN_9097; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9681 = 3'h1 == state ? dirty_1_176 : _GEN_9098; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9682 = 3'h1 == state ? dirty_1_177 : _GEN_9099; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9683 = 3'h1 == state ? dirty_1_178 : _GEN_9100; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9684 = 3'h1 == state ? dirty_1_179 : _GEN_9101; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9685 = 3'h1 == state ? dirty_1_180 : _GEN_9102; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9686 = 3'h1 == state ? dirty_1_181 : _GEN_9103; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9687 = 3'h1 == state ? dirty_1_182 : _GEN_9104; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9688 = 3'h1 == state ? dirty_1_183 : _GEN_9105; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9689 = 3'h1 == state ? dirty_1_184 : _GEN_9106; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9690 = 3'h1 == state ? dirty_1_185 : _GEN_9107; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9691 = 3'h1 == state ? dirty_1_186 : _GEN_9108; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9692 = 3'h1 == state ? dirty_1_187 : _GEN_9109; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9693 = 3'h1 == state ? dirty_1_188 : _GEN_9110; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9694 = 3'h1 == state ? dirty_1_189 : _GEN_9111; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9695 = 3'h1 == state ? dirty_1_190 : _GEN_9112; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9696 = 3'h1 == state ? dirty_1_191 : _GEN_9113; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9697 = 3'h1 == state ? dirty_1_192 : _GEN_9114; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9698 = 3'h1 == state ? dirty_1_193 : _GEN_9115; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9699 = 3'h1 == state ? dirty_1_194 : _GEN_9116; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9700 = 3'h1 == state ? dirty_1_195 : _GEN_9117; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9701 = 3'h1 == state ? dirty_1_196 : _GEN_9118; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9702 = 3'h1 == state ? dirty_1_197 : _GEN_9119; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9703 = 3'h1 == state ? dirty_1_198 : _GEN_9120; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9704 = 3'h1 == state ? dirty_1_199 : _GEN_9121; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9705 = 3'h1 == state ? dirty_1_200 : _GEN_9122; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9706 = 3'h1 == state ? dirty_1_201 : _GEN_9123; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9707 = 3'h1 == state ? dirty_1_202 : _GEN_9124; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9708 = 3'h1 == state ? dirty_1_203 : _GEN_9125; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9709 = 3'h1 == state ? dirty_1_204 : _GEN_9126; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9710 = 3'h1 == state ? dirty_1_205 : _GEN_9127; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9711 = 3'h1 == state ? dirty_1_206 : _GEN_9128; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9712 = 3'h1 == state ? dirty_1_207 : _GEN_9129; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9713 = 3'h1 == state ? dirty_1_208 : _GEN_9130; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9714 = 3'h1 == state ? dirty_1_209 : _GEN_9131; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9715 = 3'h1 == state ? dirty_1_210 : _GEN_9132; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9716 = 3'h1 == state ? dirty_1_211 : _GEN_9133; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9717 = 3'h1 == state ? dirty_1_212 : _GEN_9134; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9718 = 3'h1 == state ? dirty_1_213 : _GEN_9135; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9719 = 3'h1 == state ? dirty_1_214 : _GEN_9136; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9720 = 3'h1 == state ? dirty_1_215 : _GEN_9137; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9721 = 3'h1 == state ? dirty_1_216 : _GEN_9138; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9722 = 3'h1 == state ? dirty_1_217 : _GEN_9139; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9723 = 3'h1 == state ? dirty_1_218 : _GEN_9140; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9724 = 3'h1 == state ? dirty_1_219 : _GEN_9141; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9725 = 3'h1 == state ? dirty_1_220 : _GEN_9142; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9726 = 3'h1 == state ? dirty_1_221 : _GEN_9143; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9727 = 3'h1 == state ? dirty_1_222 : _GEN_9144; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9728 = 3'h1 == state ? dirty_1_223 : _GEN_9145; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9729 = 3'h1 == state ? dirty_1_224 : _GEN_9146; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9730 = 3'h1 == state ? dirty_1_225 : _GEN_9147; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9731 = 3'h1 == state ? dirty_1_226 : _GEN_9148; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9732 = 3'h1 == state ? dirty_1_227 : _GEN_9149; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9733 = 3'h1 == state ? dirty_1_228 : _GEN_9150; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9734 = 3'h1 == state ? dirty_1_229 : _GEN_9151; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9735 = 3'h1 == state ? dirty_1_230 : _GEN_9152; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9736 = 3'h1 == state ? dirty_1_231 : _GEN_9153; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9737 = 3'h1 == state ? dirty_1_232 : _GEN_9154; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9738 = 3'h1 == state ? dirty_1_233 : _GEN_9155; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9739 = 3'h1 == state ? dirty_1_234 : _GEN_9156; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9740 = 3'h1 == state ? dirty_1_235 : _GEN_9157; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9741 = 3'h1 == state ? dirty_1_236 : _GEN_9158; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9742 = 3'h1 == state ? dirty_1_237 : _GEN_9159; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9743 = 3'h1 == state ? dirty_1_238 : _GEN_9160; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9744 = 3'h1 == state ? dirty_1_239 : _GEN_9161; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9745 = 3'h1 == state ? dirty_1_240 : _GEN_9162; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9746 = 3'h1 == state ? dirty_1_241 : _GEN_9163; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9747 = 3'h1 == state ? dirty_1_242 : _GEN_9164; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9748 = 3'h1 == state ? dirty_1_243 : _GEN_9165; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9749 = 3'h1 == state ? dirty_1_244 : _GEN_9166; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9750 = 3'h1 == state ? dirty_1_245 : _GEN_9167; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9751 = 3'h1 == state ? dirty_1_246 : _GEN_9168; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9752 = 3'h1 == state ? dirty_1_247 : _GEN_9169; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9753 = 3'h1 == state ? dirty_1_248 : _GEN_9170; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9754 = 3'h1 == state ? dirty_1_249 : _GEN_9171; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9755 = 3'h1 == state ? dirty_1_250 : _GEN_9172; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9756 = 3'h1 == state ? dirty_1_251 : _GEN_9173; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9757 = 3'h1 == state ? dirty_1_252 : _GEN_9174; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9758 = 3'h1 == state ? dirty_1_253 : _GEN_9175; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9759 = 3'h1 == state ? dirty_1_254 : _GEN_9176; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9760 = 3'h1 == state ? dirty_1_255 : _GEN_9177; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9761 = 3'h1 == state ? 1'h0 : _GEN_9178; // @[dcache.scala 183:18 144:25]
  wire  _GEN_9762 = 3'h1 == state ? 1'h0 : _GEN_9179; // @[dcache.scala 183:18 144:25]
  wire [20:0] _GEN_9763 = 3'h1 == state ? 21'h0 : _GEN_9180; // @[dcache.scala 183:18 143:25]
  wire [20:0] _GEN_9764 = 3'h1 == state ? 21'h0 : _GEN_9181; // @[dcache.scala 183:18 143:25]
  wire [21:0] _GEN_9765 = 3'h1 == state ? 22'h0 : _GEN_9185; // @[dcache.scala 183:18 98:21]
  wire [7:0] tagv_0_addra = 3'h0 == state ? _GEN_15 : _GEN_9218; // @[dcache.scala 183:18]
  wire [31:0] _GEN_9807 = 3'h0 == state ? 32'h0 : _GEN_9233; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9808 = 3'h0 == state ? 32'h0 : _GEN_9234; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9809 = 3'h0 == state ? 32'h0 : _GEN_9235; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9810 = 3'h0 == state ? 32'h0 : _GEN_9236; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9811 = 3'h0 == state ? 32'h0 : _GEN_9237; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9812 = 3'h0 == state ? 32'h0 : _GEN_9238; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9813 = 3'h0 == state ? 32'h0 : _GEN_9239; // @[dcache.scala 183:18 149:33]
  wire [31:0] _GEN_9814 = 3'h0 == state ? 32'h0 : _GEN_9240; // @[dcache.scala 183:18 149:33]
  wire [3:0] _GEN_9815 = 3'h0 == state ? 4'h0 : _GEN_9241; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9816 = 3'h0 == state ? 4'h0 : _GEN_9242; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9817 = 3'h0 == state ? 4'h0 : _GEN_9243; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9818 = 3'h0 == state ? 4'h0 : _GEN_9244; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9819 = 3'h0 == state ? 4'h0 : _GEN_9245; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9820 = 3'h0 == state ? 4'h0 : _GEN_9246; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9821 = 3'h0 == state ? 4'h0 : _GEN_9247; // @[dcache.scala 183:18 150:33]
  wire [3:0] _GEN_9822 = 3'h0 == state ? 4'h0 : _GEN_9248; // @[dcache.scala 183:18 150:33]
  wire  _GEN_9823 = 3'h0 == state ? dirty_0_0 : _GEN_9249; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9824 = 3'h0 == state ? dirty_0_1 : _GEN_9250; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9825 = 3'h0 == state ? dirty_0_2 : _GEN_9251; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9826 = 3'h0 == state ? dirty_0_3 : _GEN_9252; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9827 = 3'h0 == state ? dirty_0_4 : _GEN_9253; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9828 = 3'h0 == state ? dirty_0_5 : _GEN_9254; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9829 = 3'h0 == state ? dirty_0_6 : _GEN_9255; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9830 = 3'h0 == state ? dirty_0_7 : _GEN_9256; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9831 = 3'h0 == state ? dirty_0_8 : _GEN_9257; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9832 = 3'h0 == state ? dirty_0_9 : _GEN_9258; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9833 = 3'h0 == state ? dirty_0_10 : _GEN_9259; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9834 = 3'h0 == state ? dirty_0_11 : _GEN_9260; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9835 = 3'h0 == state ? dirty_0_12 : _GEN_9261; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9836 = 3'h0 == state ? dirty_0_13 : _GEN_9262; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9837 = 3'h0 == state ? dirty_0_14 : _GEN_9263; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9838 = 3'h0 == state ? dirty_0_15 : _GEN_9264; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9839 = 3'h0 == state ? dirty_0_16 : _GEN_9265; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9840 = 3'h0 == state ? dirty_0_17 : _GEN_9266; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9841 = 3'h0 == state ? dirty_0_18 : _GEN_9267; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9842 = 3'h0 == state ? dirty_0_19 : _GEN_9268; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9843 = 3'h0 == state ? dirty_0_20 : _GEN_9269; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9844 = 3'h0 == state ? dirty_0_21 : _GEN_9270; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9845 = 3'h0 == state ? dirty_0_22 : _GEN_9271; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9846 = 3'h0 == state ? dirty_0_23 : _GEN_9272; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9847 = 3'h0 == state ? dirty_0_24 : _GEN_9273; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9848 = 3'h0 == state ? dirty_0_25 : _GEN_9274; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9849 = 3'h0 == state ? dirty_0_26 : _GEN_9275; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9850 = 3'h0 == state ? dirty_0_27 : _GEN_9276; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9851 = 3'h0 == state ? dirty_0_28 : _GEN_9277; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9852 = 3'h0 == state ? dirty_0_29 : _GEN_9278; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9853 = 3'h0 == state ? dirty_0_30 : _GEN_9279; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9854 = 3'h0 == state ? dirty_0_31 : _GEN_9280; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9855 = 3'h0 == state ? dirty_0_32 : _GEN_9281; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9856 = 3'h0 == state ? dirty_0_33 : _GEN_9282; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9857 = 3'h0 == state ? dirty_0_34 : _GEN_9283; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9858 = 3'h0 == state ? dirty_0_35 : _GEN_9284; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9859 = 3'h0 == state ? dirty_0_36 : _GEN_9285; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9860 = 3'h0 == state ? dirty_0_37 : _GEN_9286; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9861 = 3'h0 == state ? dirty_0_38 : _GEN_9287; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9862 = 3'h0 == state ? dirty_0_39 : _GEN_9288; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9863 = 3'h0 == state ? dirty_0_40 : _GEN_9289; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9864 = 3'h0 == state ? dirty_0_41 : _GEN_9290; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9865 = 3'h0 == state ? dirty_0_42 : _GEN_9291; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9866 = 3'h0 == state ? dirty_0_43 : _GEN_9292; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9867 = 3'h0 == state ? dirty_0_44 : _GEN_9293; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9868 = 3'h0 == state ? dirty_0_45 : _GEN_9294; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9869 = 3'h0 == state ? dirty_0_46 : _GEN_9295; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9870 = 3'h0 == state ? dirty_0_47 : _GEN_9296; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9871 = 3'h0 == state ? dirty_0_48 : _GEN_9297; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9872 = 3'h0 == state ? dirty_0_49 : _GEN_9298; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9873 = 3'h0 == state ? dirty_0_50 : _GEN_9299; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9874 = 3'h0 == state ? dirty_0_51 : _GEN_9300; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9875 = 3'h0 == state ? dirty_0_52 : _GEN_9301; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9876 = 3'h0 == state ? dirty_0_53 : _GEN_9302; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9877 = 3'h0 == state ? dirty_0_54 : _GEN_9303; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9878 = 3'h0 == state ? dirty_0_55 : _GEN_9304; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9879 = 3'h0 == state ? dirty_0_56 : _GEN_9305; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9880 = 3'h0 == state ? dirty_0_57 : _GEN_9306; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9881 = 3'h0 == state ? dirty_0_58 : _GEN_9307; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9882 = 3'h0 == state ? dirty_0_59 : _GEN_9308; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9883 = 3'h0 == state ? dirty_0_60 : _GEN_9309; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9884 = 3'h0 == state ? dirty_0_61 : _GEN_9310; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9885 = 3'h0 == state ? dirty_0_62 : _GEN_9311; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9886 = 3'h0 == state ? dirty_0_63 : _GEN_9312; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9887 = 3'h0 == state ? dirty_0_64 : _GEN_9313; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9888 = 3'h0 == state ? dirty_0_65 : _GEN_9314; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9889 = 3'h0 == state ? dirty_0_66 : _GEN_9315; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9890 = 3'h0 == state ? dirty_0_67 : _GEN_9316; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9891 = 3'h0 == state ? dirty_0_68 : _GEN_9317; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9892 = 3'h0 == state ? dirty_0_69 : _GEN_9318; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9893 = 3'h0 == state ? dirty_0_70 : _GEN_9319; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9894 = 3'h0 == state ? dirty_0_71 : _GEN_9320; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9895 = 3'h0 == state ? dirty_0_72 : _GEN_9321; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9896 = 3'h0 == state ? dirty_0_73 : _GEN_9322; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9897 = 3'h0 == state ? dirty_0_74 : _GEN_9323; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9898 = 3'h0 == state ? dirty_0_75 : _GEN_9324; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9899 = 3'h0 == state ? dirty_0_76 : _GEN_9325; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9900 = 3'h0 == state ? dirty_0_77 : _GEN_9326; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9901 = 3'h0 == state ? dirty_0_78 : _GEN_9327; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9902 = 3'h0 == state ? dirty_0_79 : _GEN_9328; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9903 = 3'h0 == state ? dirty_0_80 : _GEN_9329; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9904 = 3'h0 == state ? dirty_0_81 : _GEN_9330; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9905 = 3'h0 == state ? dirty_0_82 : _GEN_9331; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9906 = 3'h0 == state ? dirty_0_83 : _GEN_9332; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9907 = 3'h0 == state ? dirty_0_84 : _GEN_9333; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9908 = 3'h0 == state ? dirty_0_85 : _GEN_9334; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9909 = 3'h0 == state ? dirty_0_86 : _GEN_9335; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9910 = 3'h0 == state ? dirty_0_87 : _GEN_9336; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9911 = 3'h0 == state ? dirty_0_88 : _GEN_9337; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9912 = 3'h0 == state ? dirty_0_89 : _GEN_9338; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9913 = 3'h0 == state ? dirty_0_90 : _GEN_9339; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9914 = 3'h0 == state ? dirty_0_91 : _GEN_9340; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9915 = 3'h0 == state ? dirty_0_92 : _GEN_9341; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9916 = 3'h0 == state ? dirty_0_93 : _GEN_9342; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9917 = 3'h0 == state ? dirty_0_94 : _GEN_9343; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9918 = 3'h0 == state ? dirty_0_95 : _GEN_9344; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9919 = 3'h0 == state ? dirty_0_96 : _GEN_9345; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9920 = 3'h0 == state ? dirty_0_97 : _GEN_9346; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9921 = 3'h0 == state ? dirty_0_98 : _GEN_9347; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9922 = 3'h0 == state ? dirty_0_99 : _GEN_9348; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9923 = 3'h0 == state ? dirty_0_100 : _GEN_9349; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9924 = 3'h0 == state ? dirty_0_101 : _GEN_9350; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9925 = 3'h0 == state ? dirty_0_102 : _GEN_9351; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9926 = 3'h0 == state ? dirty_0_103 : _GEN_9352; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9927 = 3'h0 == state ? dirty_0_104 : _GEN_9353; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9928 = 3'h0 == state ? dirty_0_105 : _GEN_9354; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9929 = 3'h0 == state ? dirty_0_106 : _GEN_9355; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9930 = 3'h0 == state ? dirty_0_107 : _GEN_9356; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9931 = 3'h0 == state ? dirty_0_108 : _GEN_9357; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9932 = 3'h0 == state ? dirty_0_109 : _GEN_9358; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9933 = 3'h0 == state ? dirty_0_110 : _GEN_9359; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9934 = 3'h0 == state ? dirty_0_111 : _GEN_9360; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9935 = 3'h0 == state ? dirty_0_112 : _GEN_9361; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9936 = 3'h0 == state ? dirty_0_113 : _GEN_9362; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9937 = 3'h0 == state ? dirty_0_114 : _GEN_9363; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9938 = 3'h0 == state ? dirty_0_115 : _GEN_9364; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9939 = 3'h0 == state ? dirty_0_116 : _GEN_9365; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9940 = 3'h0 == state ? dirty_0_117 : _GEN_9366; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9941 = 3'h0 == state ? dirty_0_118 : _GEN_9367; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9942 = 3'h0 == state ? dirty_0_119 : _GEN_9368; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9943 = 3'h0 == state ? dirty_0_120 : _GEN_9369; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9944 = 3'h0 == state ? dirty_0_121 : _GEN_9370; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9945 = 3'h0 == state ? dirty_0_122 : _GEN_9371; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9946 = 3'h0 == state ? dirty_0_123 : _GEN_9372; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9947 = 3'h0 == state ? dirty_0_124 : _GEN_9373; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9948 = 3'h0 == state ? dirty_0_125 : _GEN_9374; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9949 = 3'h0 == state ? dirty_0_126 : _GEN_9375; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9950 = 3'h0 == state ? dirty_0_127 : _GEN_9376; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9951 = 3'h0 == state ? dirty_0_128 : _GEN_9377; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9952 = 3'h0 == state ? dirty_0_129 : _GEN_9378; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9953 = 3'h0 == state ? dirty_0_130 : _GEN_9379; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9954 = 3'h0 == state ? dirty_0_131 : _GEN_9380; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9955 = 3'h0 == state ? dirty_0_132 : _GEN_9381; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9956 = 3'h0 == state ? dirty_0_133 : _GEN_9382; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9957 = 3'h0 == state ? dirty_0_134 : _GEN_9383; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9958 = 3'h0 == state ? dirty_0_135 : _GEN_9384; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9959 = 3'h0 == state ? dirty_0_136 : _GEN_9385; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9960 = 3'h0 == state ? dirty_0_137 : _GEN_9386; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9961 = 3'h0 == state ? dirty_0_138 : _GEN_9387; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9962 = 3'h0 == state ? dirty_0_139 : _GEN_9388; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9963 = 3'h0 == state ? dirty_0_140 : _GEN_9389; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9964 = 3'h0 == state ? dirty_0_141 : _GEN_9390; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9965 = 3'h0 == state ? dirty_0_142 : _GEN_9391; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9966 = 3'h0 == state ? dirty_0_143 : _GEN_9392; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9967 = 3'h0 == state ? dirty_0_144 : _GEN_9393; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9968 = 3'h0 == state ? dirty_0_145 : _GEN_9394; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9969 = 3'h0 == state ? dirty_0_146 : _GEN_9395; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9970 = 3'h0 == state ? dirty_0_147 : _GEN_9396; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9971 = 3'h0 == state ? dirty_0_148 : _GEN_9397; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9972 = 3'h0 == state ? dirty_0_149 : _GEN_9398; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9973 = 3'h0 == state ? dirty_0_150 : _GEN_9399; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9974 = 3'h0 == state ? dirty_0_151 : _GEN_9400; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9975 = 3'h0 == state ? dirty_0_152 : _GEN_9401; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9976 = 3'h0 == state ? dirty_0_153 : _GEN_9402; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9977 = 3'h0 == state ? dirty_0_154 : _GEN_9403; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9978 = 3'h0 == state ? dirty_0_155 : _GEN_9404; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9979 = 3'h0 == state ? dirty_0_156 : _GEN_9405; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9980 = 3'h0 == state ? dirty_0_157 : _GEN_9406; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9981 = 3'h0 == state ? dirty_0_158 : _GEN_9407; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9982 = 3'h0 == state ? dirty_0_159 : _GEN_9408; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9983 = 3'h0 == state ? dirty_0_160 : _GEN_9409; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9984 = 3'h0 == state ? dirty_0_161 : _GEN_9410; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9985 = 3'h0 == state ? dirty_0_162 : _GEN_9411; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9986 = 3'h0 == state ? dirty_0_163 : _GEN_9412; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9987 = 3'h0 == state ? dirty_0_164 : _GEN_9413; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9988 = 3'h0 == state ? dirty_0_165 : _GEN_9414; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9989 = 3'h0 == state ? dirty_0_166 : _GEN_9415; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9990 = 3'h0 == state ? dirty_0_167 : _GEN_9416; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9991 = 3'h0 == state ? dirty_0_168 : _GEN_9417; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9992 = 3'h0 == state ? dirty_0_169 : _GEN_9418; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9993 = 3'h0 == state ? dirty_0_170 : _GEN_9419; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9994 = 3'h0 == state ? dirty_0_171 : _GEN_9420; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9995 = 3'h0 == state ? dirty_0_172 : _GEN_9421; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9996 = 3'h0 == state ? dirty_0_173 : _GEN_9422; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9997 = 3'h0 == state ? dirty_0_174 : _GEN_9423; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9998 = 3'h0 == state ? dirty_0_175 : _GEN_9424; // @[dcache.scala 183:18 113:28]
  wire  _GEN_9999 = 3'h0 == state ? dirty_0_176 : _GEN_9425; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10000 = 3'h0 == state ? dirty_0_177 : _GEN_9426; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10001 = 3'h0 == state ? dirty_0_178 : _GEN_9427; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10002 = 3'h0 == state ? dirty_0_179 : _GEN_9428; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10003 = 3'h0 == state ? dirty_0_180 : _GEN_9429; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10004 = 3'h0 == state ? dirty_0_181 : _GEN_9430; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10005 = 3'h0 == state ? dirty_0_182 : _GEN_9431; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10006 = 3'h0 == state ? dirty_0_183 : _GEN_9432; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10007 = 3'h0 == state ? dirty_0_184 : _GEN_9433; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10008 = 3'h0 == state ? dirty_0_185 : _GEN_9434; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10009 = 3'h0 == state ? dirty_0_186 : _GEN_9435; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10010 = 3'h0 == state ? dirty_0_187 : _GEN_9436; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10011 = 3'h0 == state ? dirty_0_188 : _GEN_9437; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10012 = 3'h0 == state ? dirty_0_189 : _GEN_9438; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10013 = 3'h0 == state ? dirty_0_190 : _GEN_9439; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10014 = 3'h0 == state ? dirty_0_191 : _GEN_9440; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10015 = 3'h0 == state ? dirty_0_192 : _GEN_9441; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10016 = 3'h0 == state ? dirty_0_193 : _GEN_9442; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10017 = 3'h0 == state ? dirty_0_194 : _GEN_9443; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10018 = 3'h0 == state ? dirty_0_195 : _GEN_9444; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10019 = 3'h0 == state ? dirty_0_196 : _GEN_9445; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10020 = 3'h0 == state ? dirty_0_197 : _GEN_9446; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10021 = 3'h0 == state ? dirty_0_198 : _GEN_9447; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10022 = 3'h0 == state ? dirty_0_199 : _GEN_9448; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10023 = 3'h0 == state ? dirty_0_200 : _GEN_9449; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10024 = 3'h0 == state ? dirty_0_201 : _GEN_9450; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10025 = 3'h0 == state ? dirty_0_202 : _GEN_9451; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10026 = 3'h0 == state ? dirty_0_203 : _GEN_9452; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10027 = 3'h0 == state ? dirty_0_204 : _GEN_9453; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10028 = 3'h0 == state ? dirty_0_205 : _GEN_9454; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10029 = 3'h0 == state ? dirty_0_206 : _GEN_9455; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10030 = 3'h0 == state ? dirty_0_207 : _GEN_9456; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10031 = 3'h0 == state ? dirty_0_208 : _GEN_9457; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10032 = 3'h0 == state ? dirty_0_209 : _GEN_9458; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10033 = 3'h0 == state ? dirty_0_210 : _GEN_9459; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10034 = 3'h0 == state ? dirty_0_211 : _GEN_9460; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10035 = 3'h0 == state ? dirty_0_212 : _GEN_9461; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10036 = 3'h0 == state ? dirty_0_213 : _GEN_9462; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10037 = 3'h0 == state ? dirty_0_214 : _GEN_9463; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10038 = 3'h0 == state ? dirty_0_215 : _GEN_9464; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10039 = 3'h0 == state ? dirty_0_216 : _GEN_9465; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10040 = 3'h0 == state ? dirty_0_217 : _GEN_9466; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10041 = 3'h0 == state ? dirty_0_218 : _GEN_9467; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10042 = 3'h0 == state ? dirty_0_219 : _GEN_9468; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10043 = 3'h0 == state ? dirty_0_220 : _GEN_9469; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10044 = 3'h0 == state ? dirty_0_221 : _GEN_9470; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10045 = 3'h0 == state ? dirty_0_222 : _GEN_9471; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10046 = 3'h0 == state ? dirty_0_223 : _GEN_9472; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10047 = 3'h0 == state ? dirty_0_224 : _GEN_9473; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10048 = 3'h0 == state ? dirty_0_225 : _GEN_9474; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10049 = 3'h0 == state ? dirty_0_226 : _GEN_9475; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10050 = 3'h0 == state ? dirty_0_227 : _GEN_9476; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10051 = 3'h0 == state ? dirty_0_228 : _GEN_9477; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10052 = 3'h0 == state ? dirty_0_229 : _GEN_9478; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10053 = 3'h0 == state ? dirty_0_230 : _GEN_9479; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10054 = 3'h0 == state ? dirty_0_231 : _GEN_9480; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10055 = 3'h0 == state ? dirty_0_232 : _GEN_9481; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10056 = 3'h0 == state ? dirty_0_233 : _GEN_9482; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10057 = 3'h0 == state ? dirty_0_234 : _GEN_9483; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10058 = 3'h0 == state ? dirty_0_235 : _GEN_9484; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10059 = 3'h0 == state ? dirty_0_236 : _GEN_9485; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10060 = 3'h0 == state ? dirty_0_237 : _GEN_9486; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10061 = 3'h0 == state ? dirty_0_238 : _GEN_9487; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10062 = 3'h0 == state ? dirty_0_239 : _GEN_9488; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10063 = 3'h0 == state ? dirty_0_240 : _GEN_9489; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10064 = 3'h0 == state ? dirty_0_241 : _GEN_9490; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10065 = 3'h0 == state ? dirty_0_242 : _GEN_9491; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10066 = 3'h0 == state ? dirty_0_243 : _GEN_9492; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10067 = 3'h0 == state ? dirty_0_244 : _GEN_9493; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10068 = 3'h0 == state ? dirty_0_245 : _GEN_9494; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10069 = 3'h0 == state ? dirty_0_246 : _GEN_9495; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10070 = 3'h0 == state ? dirty_0_247 : _GEN_9496; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10071 = 3'h0 == state ? dirty_0_248 : _GEN_9497; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10072 = 3'h0 == state ? dirty_0_249 : _GEN_9498; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10073 = 3'h0 == state ? dirty_0_250 : _GEN_9499; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10074 = 3'h0 == state ? dirty_0_251 : _GEN_9500; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10075 = 3'h0 == state ? dirty_0_252 : _GEN_9501; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10076 = 3'h0 == state ? dirty_0_253 : _GEN_9502; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10077 = 3'h0 == state ? dirty_0_254 : _GEN_9503; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10078 = 3'h0 == state ? dirty_0_255 : _GEN_9504; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10079 = 3'h0 == state ? dirty_1_0 : _GEN_9505; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10080 = 3'h0 == state ? dirty_1_1 : _GEN_9506; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10081 = 3'h0 == state ? dirty_1_2 : _GEN_9507; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10082 = 3'h0 == state ? dirty_1_3 : _GEN_9508; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10083 = 3'h0 == state ? dirty_1_4 : _GEN_9509; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10084 = 3'h0 == state ? dirty_1_5 : _GEN_9510; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10085 = 3'h0 == state ? dirty_1_6 : _GEN_9511; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10086 = 3'h0 == state ? dirty_1_7 : _GEN_9512; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10087 = 3'h0 == state ? dirty_1_8 : _GEN_9513; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10088 = 3'h0 == state ? dirty_1_9 : _GEN_9514; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10089 = 3'h0 == state ? dirty_1_10 : _GEN_9515; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10090 = 3'h0 == state ? dirty_1_11 : _GEN_9516; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10091 = 3'h0 == state ? dirty_1_12 : _GEN_9517; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10092 = 3'h0 == state ? dirty_1_13 : _GEN_9518; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10093 = 3'h0 == state ? dirty_1_14 : _GEN_9519; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10094 = 3'h0 == state ? dirty_1_15 : _GEN_9520; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10095 = 3'h0 == state ? dirty_1_16 : _GEN_9521; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10096 = 3'h0 == state ? dirty_1_17 : _GEN_9522; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10097 = 3'h0 == state ? dirty_1_18 : _GEN_9523; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10098 = 3'h0 == state ? dirty_1_19 : _GEN_9524; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10099 = 3'h0 == state ? dirty_1_20 : _GEN_9525; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10100 = 3'h0 == state ? dirty_1_21 : _GEN_9526; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10101 = 3'h0 == state ? dirty_1_22 : _GEN_9527; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10102 = 3'h0 == state ? dirty_1_23 : _GEN_9528; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10103 = 3'h0 == state ? dirty_1_24 : _GEN_9529; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10104 = 3'h0 == state ? dirty_1_25 : _GEN_9530; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10105 = 3'h0 == state ? dirty_1_26 : _GEN_9531; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10106 = 3'h0 == state ? dirty_1_27 : _GEN_9532; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10107 = 3'h0 == state ? dirty_1_28 : _GEN_9533; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10108 = 3'h0 == state ? dirty_1_29 : _GEN_9534; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10109 = 3'h0 == state ? dirty_1_30 : _GEN_9535; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10110 = 3'h0 == state ? dirty_1_31 : _GEN_9536; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10111 = 3'h0 == state ? dirty_1_32 : _GEN_9537; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10112 = 3'h0 == state ? dirty_1_33 : _GEN_9538; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10113 = 3'h0 == state ? dirty_1_34 : _GEN_9539; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10114 = 3'h0 == state ? dirty_1_35 : _GEN_9540; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10115 = 3'h0 == state ? dirty_1_36 : _GEN_9541; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10116 = 3'h0 == state ? dirty_1_37 : _GEN_9542; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10117 = 3'h0 == state ? dirty_1_38 : _GEN_9543; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10118 = 3'h0 == state ? dirty_1_39 : _GEN_9544; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10119 = 3'h0 == state ? dirty_1_40 : _GEN_9545; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10120 = 3'h0 == state ? dirty_1_41 : _GEN_9546; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10121 = 3'h0 == state ? dirty_1_42 : _GEN_9547; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10122 = 3'h0 == state ? dirty_1_43 : _GEN_9548; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10123 = 3'h0 == state ? dirty_1_44 : _GEN_9549; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10124 = 3'h0 == state ? dirty_1_45 : _GEN_9550; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10125 = 3'h0 == state ? dirty_1_46 : _GEN_9551; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10126 = 3'h0 == state ? dirty_1_47 : _GEN_9552; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10127 = 3'h0 == state ? dirty_1_48 : _GEN_9553; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10128 = 3'h0 == state ? dirty_1_49 : _GEN_9554; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10129 = 3'h0 == state ? dirty_1_50 : _GEN_9555; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10130 = 3'h0 == state ? dirty_1_51 : _GEN_9556; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10131 = 3'h0 == state ? dirty_1_52 : _GEN_9557; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10132 = 3'h0 == state ? dirty_1_53 : _GEN_9558; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10133 = 3'h0 == state ? dirty_1_54 : _GEN_9559; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10134 = 3'h0 == state ? dirty_1_55 : _GEN_9560; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10135 = 3'h0 == state ? dirty_1_56 : _GEN_9561; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10136 = 3'h0 == state ? dirty_1_57 : _GEN_9562; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10137 = 3'h0 == state ? dirty_1_58 : _GEN_9563; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10138 = 3'h0 == state ? dirty_1_59 : _GEN_9564; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10139 = 3'h0 == state ? dirty_1_60 : _GEN_9565; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10140 = 3'h0 == state ? dirty_1_61 : _GEN_9566; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10141 = 3'h0 == state ? dirty_1_62 : _GEN_9567; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10142 = 3'h0 == state ? dirty_1_63 : _GEN_9568; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10143 = 3'h0 == state ? dirty_1_64 : _GEN_9569; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10144 = 3'h0 == state ? dirty_1_65 : _GEN_9570; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10145 = 3'h0 == state ? dirty_1_66 : _GEN_9571; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10146 = 3'h0 == state ? dirty_1_67 : _GEN_9572; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10147 = 3'h0 == state ? dirty_1_68 : _GEN_9573; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10148 = 3'h0 == state ? dirty_1_69 : _GEN_9574; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10149 = 3'h0 == state ? dirty_1_70 : _GEN_9575; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10150 = 3'h0 == state ? dirty_1_71 : _GEN_9576; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10151 = 3'h0 == state ? dirty_1_72 : _GEN_9577; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10152 = 3'h0 == state ? dirty_1_73 : _GEN_9578; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10153 = 3'h0 == state ? dirty_1_74 : _GEN_9579; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10154 = 3'h0 == state ? dirty_1_75 : _GEN_9580; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10155 = 3'h0 == state ? dirty_1_76 : _GEN_9581; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10156 = 3'h0 == state ? dirty_1_77 : _GEN_9582; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10157 = 3'h0 == state ? dirty_1_78 : _GEN_9583; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10158 = 3'h0 == state ? dirty_1_79 : _GEN_9584; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10159 = 3'h0 == state ? dirty_1_80 : _GEN_9585; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10160 = 3'h0 == state ? dirty_1_81 : _GEN_9586; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10161 = 3'h0 == state ? dirty_1_82 : _GEN_9587; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10162 = 3'h0 == state ? dirty_1_83 : _GEN_9588; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10163 = 3'h0 == state ? dirty_1_84 : _GEN_9589; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10164 = 3'h0 == state ? dirty_1_85 : _GEN_9590; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10165 = 3'h0 == state ? dirty_1_86 : _GEN_9591; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10166 = 3'h0 == state ? dirty_1_87 : _GEN_9592; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10167 = 3'h0 == state ? dirty_1_88 : _GEN_9593; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10168 = 3'h0 == state ? dirty_1_89 : _GEN_9594; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10169 = 3'h0 == state ? dirty_1_90 : _GEN_9595; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10170 = 3'h0 == state ? dirty_1_91 : _GEN_9596; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10171 = 3'h0 == state ? dirty_1_92 : _GEN_9597; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10172 = 3'h0 == state ? dirty_1_93 : _GEN_9598; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10173 = 3'h0 == state ? dirty_1_94 : _GEN_9599; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10174 = 3'h0 == state ? dirty_1_95 : _GEN_9600; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10175 = 3'h0 == state ? dirty_1_96 : _GEN_9601; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10176 = 3'h0 == state ? dirty_1_97 : _GEN_9602; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10177 = 3'h0 == state ? dirty_1_98 : _GEN_9603; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10178 = 3'h0 == state ? dirty_1_99 : _GEN_9604; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10179 = 3'h0 == state ? dirty_1_100 : _GEN_9605; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10180 = 3'h0 == state ? dirty_1_101 : _GEN_9606; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10181 = 3'h0 == state ? dirty_1_102 : _GEN_9607; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10182 = 3'h0 == state ? dirty_1_103 : _GEN_9608; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10183 = 3'h0 == state ? dirty_1_104 : _GEN_9609; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10184 = 3'h0 == state ? dirty_1_105 : _GEN_9610; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10185 = 3'h0 == state ? dirty_1_106 : _GEN_9611; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10186 = 3'h0 == state ? dirty_1_107 : _GEN_9612; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10187 = 3'h0 == state ? dirty_1_108 : _GEN_9613; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10188 = 3'h0 == state ? dirty_1_109 : _GEN_9614; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10189 = 3'h0 == state ? dirty_1_110 : _GEN_9615; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10190 = 3'h0 == state ? dirty_1_111 : _GEN_9616; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10191 = 3'h0 == state ? dirty_1_112 : _GEN_9617; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10192 = 3'h0 == state ? dirty_1_113 : _GEN_9618; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10193 = 3'h0 == state ? dirty_1_114 : _GEN_9619; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10194 = 3'h0 == state ? dirty_1_115 : _GEN_9620; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10195 = 3'h0 == state ? dirty_1_116 : _GEN_9621; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10196 = 3'h0 == state ? dirty_1_117 : _GEN_9622; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10197 = 3'h0 == state ? dirty_1_118 : _GEN_9623; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10198 = 3'h0 == state ? dirty_1_119 : _GEN_9624; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10199 = 3'h0 == state ? dirty_1_120 : _GEN_9625; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10200 = 3'h0 == state ? dirty_1_121 : _GEN_9626; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10201 = 3'h0 == state ? dirty_1_122 : _GEN_9627; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10202 = 3'h0 == state ? dirty_1_123 : _GEN_9628; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10203 = 3'h0 == state ? dirty_1_124 : _GEN_9629; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10204 = 3'h0 == state ? dirty_1_125 : _GEN_9630; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10205 = 3'h0 == state ? dirty_1_126 : _GEN_9631; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10206 = 3'h0 == state ? dirty_1_127 : _GEN_9632; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10207 = 3'h0 == state ? dirty_1_128 : _GEN_9633; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10208 = 3'h0 == state ? dirty_1_129 : _GEN_9634; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10209 = 3'h0 == state ? dirty_1_130 : _GEN_9635; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10210 = 3'h0 == state ? dirty_1_131 : _GEN_9636; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10211 = 3'h0 == state ? dirty_1_132 : _GEN_9637; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10212 = 3'h0 == state ? dirty_1_133 : _GEN_9638; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10213 = 3'h0 == state ? dirty_1_134 : _GEN_9639; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10214 = 3'h0 == state ? dirty_1_135 : _GEN_9640; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10215 = 3'h0 == state ? dirty_1_136 : _GEN_9641; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10216 = 3'h0 == state ? dirty_1_137 : _GEN_9642; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10217 = 3'h0 == state ? dirty_1_138 : _GEN_9643; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10218 = 3'h0 == state ? dirty_1_139 : _GEN_9644; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10219 = 3'h0 == state ? dirty_1_140 : _GEN_9645; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10220 = 3'h0 == state ? dirty_1_141 : _GEN_9646; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10221 = 3'h0 == state ? dirty_1_142 : _GEN_9647; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10222 = 3'h0 == state ? dirty_1_143 : _GEN_9648; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10223 = 3'h0 == state ? dirty_1_144 : _GEN_9649; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10224 = 3'h0 == state ? dirty_1_145 : _GEN_9650; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10225 = 3'h0 == state ? dirty_1_146 : _GEN_9651; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10226 = 3'h0 == state ? dirty_1_147 : _GEN_9652; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10227 = 3'h0 == state ? dirty_1_148 : _GEN_9653; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10228 = 3'h0 == state ? dirty_1_149 : _GEN_9654; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10229 = 3'h0 == state ? dirty_1_150 : _GEN_9655; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10230 = 3'h0 == state ? dirty_1_151 : _GEN_9656; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10231 = 3'h0 == state ? dirty_1_152 : _GEN_9657; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10232 = 3'h0 == state ? dirty_1_153 : _GEN_9658; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10233 = 3'h0 == state ? dirty_1_154 : _GEN_9659; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10234 = 3'h0 == state ? dirty_1_155 : _GEN_9660; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10235 = 3'h0 == state ? dirty_1_156 : _GEN_9661; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10236 = 3'h0 == state ? dirty_1_157 : _GEN_9662; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10237 = 3'h0 == state ? dirty_1_158 : _GEN_9663; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10238 = 3'h0 == state ? dirty_1_159 : _GEN_9664; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10239 = 3'h0 == state ? dirty_1_160 : _GEN_9665; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10240 = 3'h0 == state ? dirty_1_161 : _GEN_9666; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10241 = 3'h0 == state ? dirty_1_162 : _GEN_9667; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10242 = 3'h0 == state ? dirty_1_163 : _GEN_9668; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10243 = 3'h0 == state ? dirty_1_164 : _GEN_9669; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10244 = 3'h0 == state ? dirty_1_165 : _GEN_9670; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10245 = 3'h0 == state ? dirty_1_166 : _GEN_9671; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10246 = 3'h0 == state ? dirty_1_167 : _GEN_9672; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10247 = 3'h0 == state ? dirty_1_168 : _GEN_9673; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10248 = 3'h0 == state ? dirty_1_169 : _GEN_9674; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10249 = 3'h0 == state ? dirty_1_170 : _GEN_9675; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10250 = 3'h0 == state ? dirty_1_171 : _GEN_9676; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10251 = 3'h0 == state ? dirty_1_172 : _GEN_9677; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10252 = 3'h0 == state ? dirty_1_173 : _GEN_9678; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10253 = 3'h0 == state ? dirty_1_174 : _GEN_9679; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10254 = 3'h0 == state ? dirty_1_175 : _GEN_9680; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10255 = 3'h0 == state ? dirty_1_176 : _GEN_9681; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10256 = 3'h0 == state ? dirty_1_177 : _GEN_9682; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10257 = 3'h0 == state ? dirty_1_178 : _GEN_9683; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10258 = 3'h0 == state ? dirty_1_179 : _GEN_9684; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10259 = 3'h0 == state ? dirty_1_180 : _GEN_9685; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10260 = 3'h0 == state ? dirty_1_181 : _GEN_9686; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10261 = 3'h0 == state ? dirty_1_182 : _GEN_9687; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10262 = 3'h0 == state ? dirty_1_183 : _GEN_9688; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10263 = 3'h0 == state ? dirty_1_184 : _GEN_9689; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10264 = 3'h0 == state ? dirty_1_185 : _GEN_9690; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10265 = 3'h0 == state ? dirty_1_186 : _GEN_9691; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10266 = 3'h0 == state ? dirty_1_187 : _GEN_9692; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10267 = 3'h0 == state ? dirty_1_188 : _GEN_9693; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10268 = 3'h0 == state ? dirty_1_189 : _GEN_9694; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10269 = 3'h0 == state ? dirty_1_190 : _GEN_9695; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10270 = 3'h0 == state ? dirty_1_191 : _GEN_9696; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10271 = 3'h0 == state ? dirty_1_192 : _GEN_9697; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10272 = 3'h0 == state ? dirty_1_193 : _GEN_9698; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10273 = 3'h0 == state ? dirty_1_194 : _GEN_9699; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10274 = 3'h0 == state ? dirty_1_195 : _GEN_9700; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10275 = 3'h0 == state ? dirty_1_196 : _GEN_9701; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10276 = 3'h0 == state ? dirty_1_197 : _GEN_9702; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10277 = 3'h0 == state ? dirty_1_198 : _GEN_9703; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10278 = 3'h0 == state ? dirty_1_199 : _GEN_9704; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10279 = 3'h0 == state ? dirty_1_200 : _GEN_9705; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10280 = 3'h0 == state ? dirty_1_201 : _GEN_9706; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10281 = 3'h0 == state ? dirty_1_202 : _GEN_9707; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10282 = 3'h0 == state ? dirty_1_203 : _GEN_9708; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10283 = 3'h0 == state ? dirty_1_204 : _GEN_9709; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10284 = 3'h0 == state ? dirty_1_205 : _GEN_9710; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10285 = 3'h0 == state ? dirty_1_206 : _GEN_9711; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10286 = 3'h0 == state ? dirty_1_207 : _GEN_9712; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10287 = 3'h0 == state ? dirty_1_208 : _GEN_9713; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10288 = 3'h0 == state ? dirty_1_209 : _GEN_9714; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10289 = 3'h0 == state ? dirty_1_210 : _GEN_9715; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10290 = 3'h0 == state ? dirty_1_211 : _GEN_9716; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10291 = 3'h0 == state ? dirty_1_212 : _GEN_9717; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10292 = 3'h0 == state ? dirty_1_213 : _GEN_9718; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10293 = 3'h0 == state ? dirty_1_214 : _GEN_9719; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10294 = 3'h0 == state ? dirty_1_215 : _GEN_9720; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10295 = 3'h0 == state ? dirty_1_216 : _GEN_9721; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10296 = 3'h0 == state ? dirty_1_217 : _GEN_9722; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10297 = 3'h0 == state ? dirty_1_218 : _GEN_9723; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10298 = 3'h0 == state ? dirty_1_219 : _GEN_9724; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10299 = 3'h0 == state ? dirty_1_220 : _GEN_9725; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10300 = 3'h0 == state ? dirty_1_221 : _GEN_9726; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10301 = 3'h0 == state ? dirty_1_222 : _GEN_9727; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10302 = 3'h0 == state ? dirty_1_223 : _GEN_9728; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10303 = 3'h0 == state ? dirty_1_224 : _GEN_9729; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10304 = 3'h0 == state ? dirty_1_225 : _GEN_9730; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10305 = 3'h0 == state ? dirty_1_226 : _GEN_9731; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10306 = 3'h0 == state ? dirty_1_227 : _GEN_9732; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10307 = 3'h0 == state ? dirty_1_228 : _GEN_9733; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10308 = 3'h0 == state ? dirty_1_229 : _GEN_9734; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10309 = 3'h0 == state ? dirty_1_230 : _GEN_9735; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10310 = 3'h0 == state ? dirty_1_231 : _GEN_9736; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10311 = 3'h0 == state ? dirty_1_232 : _GEN_9737; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10312 = 3'h0 == state ? dirty_1_233 : _GEN_9738; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10313 = 3'h0 == state ? dirty_1_234 : _GEN_9739; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10314 = 3'h0 == state ? dirty_1_235 : _GEN_9740; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10315 = 3'h0 == state ? dirty_1_236 : _GEN_9741; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10316 = 3'h0 == state ? dirty_1_237 : _GEN_9742; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10317 = 3'h0 == state ? dirty_1_238 : _GEN_9743; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10318 = 3'h0 == state ? dirty_1_239 : _GEN_9744; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10319 = 3'h0 == state ? dirty_1_240 : _GEN_9745; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10320 = 3'h0 == state ? dirty_1_241 : _GEN_9746; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10321 = 3'h0 == state ? dirty_1_242 : _GEN_9747; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10322 = 3'h0 == state ? dirty_1_243 : _GEN_9748; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10323 = 3'h0 == state ? dirty_1_244 : _GEN_9749; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10324 = 3'h0 == state ? dirty_1_245 : _GEN_9750; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10325 = 3'h0 == state ? dirty_1_246 : _GEN_9751; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10326 = 3'h0 == state ? dirty_1_247 : _GEN_9752; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10327 = 3'h0 == state ? dirty_1_248 : _GEN_9753; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10328 = 3'h0 == state ? dirty_1_249 : _GEN_9754; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10329 = 3'h0 == state ? dirty_1_250 : _GEN_9755; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10330 = 3'h0 == state ? dirty_1_251 : _GEN_9756; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10331 = 3'h0 == state ? dirty_1_252 : _GEN_9757; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10332 = 3'h0 == state ? dirty_1_253 : _GEN_9758; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10333 = 3'h0 == state ? dirty_1_254 : _GEN_9759; // @[dcache.scala 183:18 113:28]
  wire  _GEN_10334 = 3'h0 == state ? dirty_1_255 : _GEN_9760; // @[dcache.scala 183:18 113:28]
  wire  _T_53 = hit & req_op; // @[dcache.scala 448:22]
  wire  _GEN_16590 = ~req_wline; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10341 = ~req_wline & 8'h0 == req_wset | _GEN_9823; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10342 = ~req_wline & 8'h1 == req_wset | _GEN_9824; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10343 = ~req_wline & 8'h2 == req_wset | _GEN_9825; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10344 = ~req_wline & 8'h3 == req_wset | _GEN_9826; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10345 = ~req_wline & 8'h4 == req_wset | _GEN_9827; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10346 = ~req_wline & 8'h5 == req_wset | _GEN_9828; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10347 = ~req_wline & 8'h6 == req_wset | _GEN_9829; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10348 = ~req_wline & 8'h7 == req_wset | _GEN_9830; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10349 = ~req_wline & 8'h8 == req_wset | _GEN_9831; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10350 = ~req_wline & 8'h9 == req_wset | _GEN_9832; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10351 = ~req_wline & 8'ha == req_wset | _GEN_9833; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10352 = ~req_wline & 8'hb == req_wset | _GEN_9834; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10353 = ~req_wline & 8'hc == req_wset | _GEN_9835; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10354 = ~req_wline & 8'hd == req_wset | _GEN_9836; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10355 = ~req_wline & 8'he == req_wset | _GEN_9837; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10356 = ~req_wline & 8'hf == req_wset | _GEN_9838; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10357 = ~req_wline & 8'h10 == req_wset | _GEN_9839; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10358 = ~req_wline & 8'h11 == req_wset | _GEN_9840; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10359 = ~req_wline & 8'h12 == req_wset | _GEN_9841; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10360 = ~req_wline & 8'h13 == req_wset | _GEN_9842; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10361 = ~req_wline & 8'h14 == req_wset | _GEN_9843; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10362 = ~req_wline & 8'h15 == req_wset | _GEN_9844; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10363 = ~req_wline & 8'h16 == req_wset | _GEN_9845; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10364 = ~req_wline & 8'h17 == req_wset | _GEN_9846; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10365 = ~req_wline & 8'h18 == req_wset | _GEN_9847; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10366 = ~req_wline & 8'h19 == req_wset | _GEN_9848; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10367 = ~req_wline & 8'h1a == req_wset | _GEN_9849; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10368 = ~req_wline & 8'h1b == req_wset | _GEN_9850; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10369 = ~req_wline & 8'h1c == req_wset | _GEN_9851; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10370 = ~req_wline & 8'h1d == req_wset | _GEN_9852; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10371 = ~req_wline & 8'h1e == req_wset | _GEN_9853; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10372 = ~req_wline & 8'h1f == req_wset | _GEN_9854; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10373 = ~req_wline & 8'h20 == req_wset | _GEN_9855; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10374 = ~req_wline & 8'h21 == req_wset | _GEN_9856; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10375 = ~req_wline & 8'h22 == req_wset | _GEN_9857; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10376 = ~req_wline & 8'h23 == req_wset | _GEN_9858; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10377 = ~req_wline & 8'h24 == req_wset | _GEN_9859; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10378 = ~req_wline & 8'h25 == req_wset | _GEN_9860; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10379 = ~req_wline & 8'h26 == req_wset | _GEN_9861; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10380 = ~req_wline & 8'h27 == req_wset | _GEN_9862; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10381 = ~req_wline & 8'h28 == req_wset | _GEN_9863; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10382 = ~req_wline & 8'h29 == req_wset | _GEN_9864; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10383 = ~req_wline & 8'h2a == req_wset | _GEN_9865; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10384 = ~req_wline & 8'h2b == req_wset | _GEN_9866; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10385 = ~req_wline & 8'h2c == req_wset | _GEN_9867; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10386 = ~req_wline & 8'h2d == req_wset | _GEN_9868; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10387 = ~req_wline & 8'h2e == req_wset | _GEN_9869; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10388 = ~req_wline & 8'h2f == req_wset | _GEN_9870; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10389 = ~req_wline & 8'h30 == req_wset | _GEN_9871; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10390 = ~req_wline & 8'h31 == req_wset | _GEN_9872; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10391 = ~req_wline & 8'h32 == req_wset | _GEN_9873; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10392 = ~req_wline & 8'h33 == req_wset | _GEN_9874; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10393 = ~req_wline & 8'h34 == req_wset | _GEN_9875; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10394 = ~req_wline & 8'h35 == req_wset | _GEN_9876; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10395 = ~req_wline & 8'h36 == req_wset | _GEN_9877; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10396 = ~req_wline & 8'h37 == req_wset | _GEN_9878; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10397 = ~req_wline & 8'h38 == req_wset | _GEN_9879; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10398 = ~req_wline & 8'h39 == req_wset | _GEN_9880; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10399 = ~req_wline & 8'h3a == req_wset | _GEN_9881; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10400 = ~req_wline & 8'h3b == req_wset | _GEN_9882; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10401 = ~req_wline & 8'h3c == req_wset | _GEN_9883; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10402 = ~req_wline & 8'h3d == req_wset | _GEN_9884; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10403 = ~req_wline & 8'h3e == req_wset | _GEN_9885; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10404 = ~req_wline & 8'h3f == req_wset | _GEN_9886; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10405 = ~req_wline & 8'h40 == req_wset | _GEN_9887; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10406 = ~req_wline & 8'h41 == req_wset | _GEN_9888; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10407 = ~req_wline & 8'h42 == req_wset | _GEN_9889; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10408 = ~req_wline & 8'h43 == req_wset | _GEN_9890; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10409 = ~req_wline & 8'h44 == req_wset | _GEN_9891; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10410 = ~req_wline & 8'h45 == req_wset | _GEN_9892; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10411 = ~req_wline & 8'h46 == req_wset | _GEN_9893; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10412 = ~req_wline & 8'h47 == req_wset | _GEN_9894; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10413 = ~req_wline & 8'h48 == req_wset | _GEN_9895; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10414 = ~req_wline & 8'h49 == req_wset | _GEN_9896; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10415 = ~req_wline & 8'h4a == req_wset | _GEN_9897; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10416 = ~req_wline & 8'h4b == req_wset | _GEN_9898; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10417 = ~req_wline & 8'h4c == req_wset | _GEN_9899; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10418 = ~req_wline & 8'h4d == req_wset | _GEN_9900; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10419 = ~req_wline & 8'h4e == req_wset | _GEN_9901; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10420 = ~req_wline & 8'h4f == req_wset | _GEN_9902; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10421 = ~req_wline & 8'h50 == req_wset | _GEN_9903; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10422 = ~req_wline & 8'h51 == req_wset | _GEN_9904; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10423 = ~req_wline & 8'h52 == req_wset | _GEN_9905; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10424 = ~req_wline & 8'h53 == req_wset | _GEN_9906; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10425 = ~req_wline & 8'h54 == req_wset | _GEN_9907; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10426 = ~req_wline & 8'h55 == req_wset | _GEN_9908; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10427 = ~req_wline & 8'h56 == req_wset | _GEN_9909; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10428 = ~req_wline & 8'h57 == req_wset | _GEN_9910; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10429 = ~req_wline & 8'h58 == req_wset | _GEN_9911; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10430 = ~req_wline & 8'h59 == req_wset | _GEN_9912; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10431 = ~req_wline & 8'h5a == req_wset | _GEN_9913; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10432 = ~req_wline & 8'h5b == req_wset | _GEN_9914; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10433 = ~req_wline & 8'h5c == req_wset | _GEN_9915; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10434 = ~req_wline & 8'h5d == req_wset | _GEN_9916; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10435 = ~req_wline & 8'h5e == req_wset | _GEN_9917; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10436 = ~req_wline & 8'h5f == req_wset | _GEN_9918; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10437 = ~req_wline & 8'h60 == req_wset | _GEN_9919; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10438 = ~req_wline & 8'h61 == req_wset | _GEN_9920; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10439 = ~req_wline & 8'h62 == req_wset | _GEN_9921; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10440 = ~req_wline & 8'h63 == req_wset | _GEN_9922; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10441 = ~req_wline & 8'h64 == req_wset | _GEN_9923; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10442 = ~req_wline & 8'h65 == req_wset | _GEN_9924; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10443 = ~req_wline & 8'h66 == req_wset | _GEN_9925; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10444 = ~req_wline & 8'h67 == req_wset | _GEN_9926; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10445 = ~req_wline & 8'h68 == req_wset | _GEN_9927; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10446 = ~req_wline & 8'h69 == req_wset | _GEN_9928; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10447 = ~req_wline & 8'h6a == req_wset | _GEN_9929; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10448 = ~req_wline & 8'h6b == req_wset | _GEN_9930; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10449 = ~req_wline & 8'h6c == req_wset | _GEN_9931; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10450 = ~req_wline & 8'h6d == req_wset | _GEN_9932; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10451 = ~req_wline & 8'h6e == req_wset | _GEN_9933; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10452 = ~req_wline & 8'h6f == req_wset | _GEN_9934; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10453 = ~req_wline & 8'h70 == req_wset | _GEN_9935; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10454 = ~req_wline & 8'h71 == req_wset | _GEN_9936; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10455 = ~req_wline & 8'h72 == req_wset | _GEN_9937; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10456 = ~req_wline & 8'h73 == req_wset | _GEN_9938; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10457 = ~req_wline & 8'h74 == req_wset | _GEN_9939; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10458 = ~req_wline & 8'h75 == req_wset | _GEN_9940; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10459 = ~req_wline & 8'h76 == req_wset | _GEN_9941; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10460 = ~req_wline & 8'h77 == req_wset | _GEN_9942; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10461 = ~req_wline & 8'h78 == req_wset | _GEN_9943; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10462 = ~req_wline & 8'h79 == req_wset | _GEN_9944; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10463 = ~req_wline & 8'h7a == req_wset | _GEN_9945; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10464 = ~req_wline & 8'h7b == req_wset | _GEN_9946; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10465 = ~req_wline & 8'h7c == req_wset | _GEN_9947; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10466 = ~req_wline & 8'h7d == req_wset | _GEN_9948; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10467 = ~req_wline & 8'h7e == req_wset | _GEN_9949; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10468 = ~req_wline & 8'h7f == req_wset | _GEN_9950; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10469 = ~req_wline & 8'h80 == req_wset | _GEN_9951; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10470 = ~req_wline & 8'h81 == req_wset | _GEN_9952; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10471 = ~req_wline & 8'h82 == req_wset | _GEN_9953; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10472 = ~req_wline & 8'h83 == req_wset | _GEN_9954; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10473 = ~req_wline & 8'h84 == req_wset | _GEN_9955; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10474 = ~req_wline & 8'h85 == req_wset | _GEN_9956; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10475 = ~req_wline & 8'h86 == req_wset | _GEN_9957; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10476 = ~req_wline & 8'h87 == req_wset | _GEN_9958; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10477 = ~req_wline & 8'h88 == req_wset | _GEN_9959; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10478 = ~req_wline & 8'h89 == req_wset | _GEN_9960; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10479 = ~req_wline & 8'h8a == req_wset | _GEN_9961; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10480 = ~req_wline & 8'h8b == req_wset | _GEN_9962; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10481 = ~req_wline & 8'h8c == req_wset | _GEN_9963; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10482 = ~req_wline & 8'h8d == req_wset | _GEN_9964; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10483 = ~req_wline & 8'h8e == req_wset | _GEN_9965; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10484 = ~req_wline & 8'h8f == req_wset | _GEN_9966; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10485 = ~req_wline & 8'h90 == req_wset | _GEN_9967; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10486 = ~req_wline & 8'h91 == req_wset | _GEN_9968; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10487 = ~req_wline & 8'h92 == req_wset | _GEN_9969; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10488 = ~req_wline & 8'h93 == req_wset | _GEN_9970; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10489 = ~req_wline & 8'h94 == req_wset | _GEN_9971; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10490 = ~req_wline & 8'h95 == req_wset | _GEN_9972; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10491 = ~req_wline & 8'h96 == req_wset | _GEN_9973; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10492 = ~req_wline & 8'h97 == req_wset | _GEN_9974; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10493 = ~req_wline & 8'h98 == req_wset | _GEN_9975; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10494 = ~req_wline & 8'h99 == req_wset | _GEN_9976; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10495 = ~req_wline & 8'h9a == req_wset | _GEN_9977; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10496 = ~req_wline & 8'h9b == req_wset | _GEN_9978; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10497 = ~req_wline & 8'h9c == req_wset | _GEN_9979; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10498 = ~req_wline & 8'h9d == req_wset | _GEN_9980; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10499 = ~req_wline & 8'h9e == req_wset | _GEN_9981; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10500 = ~req_wline & 8'h9f == req_wset | _GEN_9982; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10501 = ~req_wline & 8'ha0 == req_wset | _GEN_9983; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10502 = ~req_wline & 8'ha1 == req_wset | _GEN_9984; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10503 = ~req_wline & 8'ha2 == req_wset | _GEN_9985; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10504 = ~req_wline & 8'ha3 == req_wset | _GEN_9986; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10505 = ~req_wline & 8'ha4 == req_wset | _GEN_9987; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10506 = ~req_wline & 8'ha5 == req_wset | _GEN_9988; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10507 = ~req_wline & 8'ha6 == req_wset | _GEN_9989; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10508 = ~req_wline & 8'ha7 == req_wset | _GEN_9990; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10509 = ~req_wline & 8'ha8 == req_wset | _GEN_9991; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10510 = ~req_wline & 8'ha9 == req_wset | _GEN_9992; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10511 = ~req_wline & 8'haa == req_wset | _GEN_9993; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10512 = ~req_wline & 8'hab == req_wset | _GEN_9994; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10513 = ~req_wline & 8'hac == req_wset | _GEN_9995; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10514 = ~req_wline & 8'had == req_wset | _GEN_9996; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10515 = ~req_wline & 8'hae == req_wset | _GEN_9997; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10516 = ~req_wline & 8'haf == req_wset | _GEN_9998; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10517 = ~req_wline & 8'hb0 == req_wset | _GEN_9999; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10518 = ~req_wline & 8'hb1 == req_wset | _GEN_10000; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10519 = ~req_wline & 8'hb2 == req_wset | _GEN_10001; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10520 = ~req_wline & 8'hb3 == req_wset | _GEN_10002; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10521 = ~req_wline & 8'hb4 == req_wset | _GEN_10003; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10522 = ~req_wline & 8'hb5 == req_wset | _GEN_10004; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10523 = ~req_wline & 8'hb6 == req_wset | _GEN_10005; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10524 = ~req_wline & 8'hb7 == req_wset | _GEN_10006; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10525 = ~req_wline & 8'hb8 == req_wset | _GEN_10007; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10526 = ~req_wline & 8'hb9 == req_wset | _GEN_10008; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10527 = ~req_wline & 8'hba == req_wset | _GEN_10009; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10528 = ~req_wline & 8'hbb == req_wset | _GEN_10010; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10529 = ~req_wline & 8'hbc == req_wset | _GEN_10011; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10530 = ~req_wline & 8'hbd == req_wset | _GEN_10012; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10531 = ~req_wline & 8'hbe == req_wset | _GEN_10013; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10532 = ~req_wline & 8'hbf == req_wset | _GEN_10014; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10533 = ~req_wline & 8'hc0 == req_wset | _GEN_10015; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10534 = ~req_wline & 8'hc1 == req_wset | _GEN_10016; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10535 = ~req_wline & 8'hc2 == req_wset | _GEN_10017; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10536 = ~req_wline & 8'hc3 == req_wset | _GEN_10018; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10537 = ~req_wline & 8'hc4 == req_wset | _GEN_10019; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10538 = ~req_wline & 8'hc5 == req_wset | _GEN_10020; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10539 = ~req_wline & 8'hc6 == req_wset | _GEN_10021; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10540 = ~req_wline & 8'hc7 == req_wset | _GEN_10022; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10541 = ~req_wline & 8'hc8 == req_wset | _GEN_10023; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10542 = ~req_wline & 8'hc9 == req_wset | _GEN_10024; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10543 = ~req_wline & 8'hca == req_wset | _GEN_10025; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10544 = ~req_wline & 8'hcb == req_wset | _GEN_10026; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10545 = ~req_wline & 8'hcc == req_wset | _GEN_10027; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10546 = ~req_wline & 8'hcd == req_wset | _GEN_10028; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10547 = ~req_wline & 8'hce == req_wset | _GEN_10029; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10548 = ~req_wline & 8'hcf == req_wset | _GEN_10030; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10549 = ~req_wline & 8'hd0 == req_wset | _GEN_10031; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10550 = ~req_wline & 8'hd1 == req_wset | _GEN_10032; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10551 = ~req_wline & 8'hd2 == req_wset | _GEN_10033; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10552 = ~req_wline & 8'hd3 == req_wset | _GEN_10034; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10553 = ~req_wline & 8'hd4 == req_wset | _GEN_10035; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10554 = ~req_wline & 8'hd5 == req_wset | _GEN_10036; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10555 = ~req_wline & 8'hd6 == req_wset | _GEN_10037; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10556 = ~req_wline & 8'hd7 == req_wset | _GEN_10038; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10557 = ~req_wline & 8'hd8 == req_wset | _GEN_10039; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10558 = ~req_wline & 8'hd9 == req_wset | _GEN_10040; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10559 = ~req_wline & 8'hda == req_wset | _GEN_10041; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10560 = ~req_wline & 8'hdb == req_wset | _GEN_10042; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10561 = ~req_wline & 8'hdc == req_wset | _GEN_10043; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10562 = ~req_wline & 8'hdd == req_wset | _GEN_10044; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10563 = ~req_wline & 8'hde == req_wset | _GEN_10045; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10564 = ~req_wline & 8'hdf == req_wset | _GEN_10046; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10565 = ~req_wline & 8'he0 == req_wset | _GEN_10047; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10566 = ~req_wline & 8'he1 == req_wset | _GEN_10048; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10567 = ~req_wline & 8'he2 == req_wset | _GEN_10049; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10568 = ~req_wline & 8'he3 == req_wset | _GEN_10050; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10569 = ~req_wline & 8'he4 == req_wset | _GEN_10051; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10570 = ~req_wline & 8'he5 == req_wset | _GEN_10052; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10571 = ~req_wline & 8'he6 == req_wset | _GEN_10053; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10572 = ~req_wline & 8'he7 == req_wset | _GEN_10054; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10573 = ~req_wline & 8'he8 == req_wset | _GEN_10055; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10574 = ~req_wline & 8'he9 == req_wset | _GEN_10056; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10575 = ~req_wline & 8'hea == req_wset | _GEN_10057; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10576 = ~req_wline & 8'heb == req_wset | _GEN_10058; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10577 = ~req_wline & 8'hec == req_wset | _GEN_10059; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10578 = ~req_wline & 8'hed == req_wset | _GEN_10060; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10579 = ~req_wline & 8'hee == req_wset | _GEN_10061; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10580 = ~req_wline & 8'hef == req_wset | _GEN_10062; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10581 = ~req_wline & 8'hf0 == req_wset | _GEN_10063; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10582 = ~req_wline & 8'hf1 == req_wset | _GEN_10064; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10583 = ~req_wline & 8'hf2 == req_wset | _GEN_10065; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10584 = ~req_wline & 8'hf3 == req_wset | _GEN_10066; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10585 = ~req_wline & 8'hf4 == req_wset | _GEN_10067; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10586 = ~req_wline & 8'hf5 == req_wset | _GEN_10068; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10587 = ~req_wline & 8'hf6 == req_wset | _GEN_10069; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10588 = ~req_wline & 8'hf7 == req_wset | _GEN_10070; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10589 = ~req_wline & 8'hf8 == req_wset | _GEN_10071; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10590 = ~req_wline & 8'hf9 == req_wset | _GEN_10072; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10591 = ~req_wline & 8'hfa == req_wset | _GEN_10073; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10592 = ~req_wline & 8'hfb == req_wset | _GEN_10074; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10593 = ~req_wline & 8'hfc == req_wset | _GEN_10075; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10594 = ~req_wline & 8'hfd == req_wset | _GEN_10076; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10595 = ~req_wline & 8'hfe == req_wset | _GEN_10077; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10596 = ~req_wline & 8'hff == req_wset | _GEN_10078; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10597 = req_wline & 8'h0 == req_wset | _GEN_10079; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10598 = req_wline & 8'h1 == req_wset | _GEN_10080; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10599 = req_wline & 8'h2 == req_wset | _GEN_10081; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10600 = req_wline & 8'h3 == req_wset | _GEN_10082; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10601 = req_wline & 8'h4 == req_wset | _GEN_10083; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10602 = req_wline & 8'h5 == req_wset | _GEN_10084; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10603 = req_wline & 8'h6 == req_wset | _GEN_10085; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10604 = req_wline & 8'h7 == req_wset | _GEN_10086; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10605 = req_wline & 8'h8 == req_wset | _GEN_10087; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10606 = req_wline & 8'h9 == req_wset | _GEN_10088; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10607 = req_wline & 8'ha == req_wset | _GEN_10089; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10608 = req_wline & 8'hb == req_wset | _GEN_10090; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10609 = req_wline & 8'hc == req_wset | _GEN_10091; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10610 = req_wline & 8'hd == req_wset | _GEN_10092; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10611 = req_wline & 8'he == req_wset | _GEN_10093; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10612 = req_wline & 8'hf == req_wset | _GEN_10094; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10613 = req_wline & 8'h10 == req_wset | _GEN_10095; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10614 = req_wline & 8'h11 == req_wset | _GEN_10096; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10615 = req_wline & 8'h12 == req_wset | _GEN_10097; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10616 = req_wline & 8'h13 == req_wset | _GEN_10098; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10617 = req_wline & 8'h14 == req_wset | _GEN_10099; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10618 = req_wline & 8'h15 == req_wset | _GEN_10100; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10619 = req_wline & 8'h16 == req_wset | _GEN_10101; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10620 = req_wline & 8'h17 == req_wset | _GEN_10102; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10621 = req_wline & 8'h18 == req_wset | _GEN_10103; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10622 = req_wline & 8'h19 == req_wset | _GEN_10104; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10623 = req_wline & 8'h1a == req_wset | _GEN_10105; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10624 = req_wline & 8'h1b == req_wset | _GEN_10106; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10625 = req_wline & 8'h1c == req_wset | _GEN_10107; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10626 = req_wline & 8'h1d == req_wset | _GEN_10108; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10627 = req_wline & 8'h1e == req_wset | _GEN_10109; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10628 = req_wline & 8'h1f == req_wset | _GEN_10110; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10629 = req_wline & 8'h20 == req_wset | _GEN_10111; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10630 = req_wline & 8'h21 == req_wset | _GEN_10112; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10631 = req_wline & 8'h22 == req_wset | _GEN_10113; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10632 = req_wline & 8'h23 == req_wset | _GEN_10114; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10633 = req_wline & 8'h24 == req_wset | _GEN_10115; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10634 = req_wline & 8'h25 == req_wset | _GEN_10116; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10635 = req_wline & 8'h26 == req_wset | _GEN_10117; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10636 = req_wline & 8'h27 == req_wset | _GEN_10118; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10637 = req_wline & 8'h28 == req_wset | _GEN_10119; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10638 = req_wline & 8'h29 == req_wset | _GEN_10120; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10639 = req_wline & 8'h2a == req_wset | _GEN_10121; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10640 = req_wline & 8'h2b == req_wset | _GEN_10122; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10641 = req_wline & 8'h2c == req_wset | _GEN_10123; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10642 = req_wline & 8'h2d == req_wset | _GEN_10124; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10643 = req_wline & 8'h2e == req_wset | _GEN_10125; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10644 = req_wline & 8'h2f == req_wset | _GEN_10126; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10645 = req_wline & 8'h30 == req_wset | _GEN_10127; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10646 = req_wline & 8'h31 == req_wset | _GEN_10128; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10647 = req_wline & 8'h32 == req_wset | _GEN_10129; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10648 = req_wline & 8'h33 == req_wset | _GEN_10130; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10649 = req_wline & 8'h34 == req_wset | _GEN_10131; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10650 = req_wline & 8'h35 == req_wset | _GEN_10132; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10651 = req_wline & 8'h36 == req_wset | _GEN_10133; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10652 = req_wline & 8'h37 == req_wset | _GEN_10134; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10653 = req_wline & 8'h38 == req_wset | _GEN_10135; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10654 = req_wline & 8'h39 == req_wset | _GEN_10136; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10655 = req_wline & 8'h3a == req_wset | _GEN_10137; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10656 = req_wline & 8'h3b == req_wset | _GEN_10138; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10657 = req_wline & 8'h3c == req_wset | _GEN_10139; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10658 = req_wline & 8'h3d == req_wset | _GEN_10140; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10659 = req_wline & 8'h3e == req_wset | _GEN_10141; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10660 = req_wline & 8'h3f == req_wset | _GEN_10142; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10661 = req_wline & 8'h40 == req_wset | _GEN_10143; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10662 = req_wline & 8'h41 == req_wset | _GEN_10144; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10663 = req_wline & 8'h42 == req_wset | _GEN_10145; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10664 = req_wline & 8'h43 == req_wset | _GEN_10146; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10665 = req_wline & 8'h44 == req_wset | _GEN_10147; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10666 = req_wline & 8'h45 == req_wset | _GEN_10148; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10667 = req_wline & 8'h46 == req_wset | _GEN_10149; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10668 = req_wline & 8'h47 == req_wset | _GEN_10150; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10669 = req_wline & 8'h48 == req_wset | _GEN_10151; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10670 = req_wline & 8'h49 == req_wset | _GEN_10152; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10671 = req_wline & 8'h4a == req_wset | _GEN_10153; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10672 = req_wline & 8'h4b == req_wset | _GEN_10154; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10673 = req_wline & 8'h4c == req_wset | _GEN_10155; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10674 = req_wline & 8'h4d == req_wset | _GEN_10156; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10675 = req_wline & 8'h4e == req_wset | _GEN_10157; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10676 = req_wline & 8'h4f == req_wset | _GEN_10158; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10677 = req_wline & 8'h50 == req_wset | _GEN_10159; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10678 = req_wline & 8'h51 == req_wset | _GEN_10160; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10679 = req_wline & 8'h52 == req_wset | _GEN_10161; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10680 = req_wline & 8'h53 == req_wset | _GEN_10162; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10681 = req_wline & 8'h54 == req_wset | _GEN_10163; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10682 = req_wline & 8'h55 == req_wset | _GEN_10164; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10683 = req_wline & 8'h56 == req_wset | _GEN_10165; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10684 = req_wline & 8'h57 == req_wset | _GEN_10166; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10685 = req_wline & 8'h58 == req_wset | _GEN_10167; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10686 = req_wline & 8'h59 == req_wset | _GEN_10168; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10687 = req_wline & 8'h5a == req_wset | _GEN_10169; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10688 = req_wline & 8'h5b == req_wset | _GEN_10170; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10689 = req_wline & 8'h5c == req_wset | _GEN_10171; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10690 = req_wline & 8'h5d == req_wset | _GEN_10172; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10691 = req_wline & 8'h5e == req_wset | _GEN_10173; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10692 = req_wline & 8'h5f == req_wset | _GEN_10174; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10693 = req_wline & 8'h60 == req_wset | _GEN_10175; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10694 = req_wline & 8'h61 == req_wset | _GEN_10176; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10695 = req_wline & 8'h62 == req_wset | _GEN_10177; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10696 = req_wline & 8'h63 == req_wset | _GEN_10178; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10697 = req_wline & 8'h64 == req_wset | _GEN_10179; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10698 = req_wline & 8'h65 == req_wset | _GEN_10180; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10699 = req_wline & 8'h66 == req_wset | _GEN_10181; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10700 = req_wline & 8'h67 == req_wset | _GEN_10182; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10701 = req_wline & 8'h68 == req_wset | _GEN_10183; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10702 = req_wline & 8'h69 == req_wset | _GEN_10184; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10703 = req_wline & 8'h6a == req_wset | _GEN_10185; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10704 = req_wline & 8'h6b == req_wset | _GEN_10186; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10705 = req_wline & 8'h6c == req_wset | _GEN_10187; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10706 = req_wline & 8'h6d == req_wset | _GEN_10188; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10707 = req_wline & 8'h6e == req_wset | _GEN_10189; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10708 = req_wline & 8'h6f == req_wset | _GEN_10190; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10709 = req_wline & 8'h70 == req_wset | _GEN_10191; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10710 = req_wline & 8'h71 == req_wset | _GEN_10192; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10711 = req_wline & 8'h72 == req_wset | _GEN_10193; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10712 = req_wline & 8'h73 == req_wset | _GEN_10194; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10713 = req_wline & 8'h74 == req_wset | _GEN_10195; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10714 = req_wline & 8'h75 == req_wset | _GEN_10196; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10715 = req_wline & 8'h76 == req_wset | _GEN_10197; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10716 = req_wline & 8'h77 == req_wset | _GEN_10198; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10717 = req_wline & 8'h78 == req_wset | _GEN_10199; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10718 = req_wline & 8'h79 == req_wset | _GEN_10200; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10719 = req_wline & 8'h7a == req_wset | _GEN_10201; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10720 = req_wline & 8'h7b == req_wset | _GEN_10202; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10721 = req_wline & 8'h7c == req_wset | _GEN_10203; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10722 = req_wline & 8'h7d == req_wset | _GEN_10204; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10723 = req_wline & 8'h7e == req_wset | _GEN_10205; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10724 = req_wline & 8'h7f == req_wset | _GEN_10206; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10725 = req_wline & 8'h80 == req_wset | _GEN_10207; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10726 = req_wline & 8'h81 == req_wset | _GEN_10208; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10727 = req_wline & 8'h82 == req_wset | _GEN_10209; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10728 = req_wline & 8'h83 == req_wset | _GEN_10210; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10729 = req_wline & 8'h84 == req_wset | _GEN_10211; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10730 = req_wline & 8'h85 == req_wset | _GEN_10212; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10731 = req_wline & 8'h86 == req_wset | _GEN_10213; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10732 = req_wline & 8'h87 == req_wset | _GEN_10214; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10733 = req_wline & 8'h88 == req_wset | _GEN_10215; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10734 = req_wline & 8'h89 == req_wset | _GEN_10216; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10735 = req_wline & 8'h8a == req_wset | _GEN_10217; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10736 = req_wline & 8'h8b == req_wset | _GEN_10218; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10737 = req_wline & 8'h8c == req_wset | _GEN_10219; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10738 = req_wline & 8'h8d == req_wset | _GEN_10220; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10739 = req_wline & 8'h8e == req_wset | _GEN_10221; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10740 = req_wline & 8'h8f == req_wset | _GEN_10222; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10741 = req_wline & 8'h90 == req_wset | _GEN_10223; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10742 = req_wline & 8'h91 == req_wset | _GEN_10224; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10743 = req_wline & 8'h92 == req_wset | _GEN_10225; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10744 = req_wline & 8'h93 == req_wset | _GEN_10226; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10745 = req_wline & 8'h94 == req_wset | _GEN_10227; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10746 = req_wline & 8'h95 == req_wset | _GEN_10228; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10747 = req_wline & 8'h96 == req_wset | _GEN_10229; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10748 = req_wline & 8'h97 == req_wset | _GEN_10230; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10749 = req_wline & 8'h98 == req_wset | _GEN_10231; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10750 = req_wline & 8'h99 == req_wset | _GEN_10232; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10751 = req_wline & 8'h9a == req_wset | _GEN_10233; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10752 = req_wline & 8'h9b == req_wset | _GEN_10234; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10753 = req_wline & 8'h9c == req_wset | _GEN_10235; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10754 = req_wline & 8'h9d == req_wset | _GEN_10236; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10755 = req_wline & 8'h9e == req_wset | _GEN_10237; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10756 = req_wline & 8'h9f == req_wset | _GEN_10238; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10757 = req_wline & 8'ha0 == req_wset | _GEN_10239; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10758 = req_wline & 8'ha1 == req_wset | _GEN_10240; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10759 = req_wline & 8'ha2 == req_wset | _GEN_10241; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10760 = req_wline & 8'ha3 == req_wset | _GEN_10242; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10761 = req_wline & 8'ha4 == req_wset | _GEN_10243; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10762 = req_wline & 8'ha5 == req_wset | _GEN_10244; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10763 = req_wline & 8'ha6 == req_wset | _GEN_10245; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10764 = req_wline & 8'ha7 == req_wset | _GEN_10246; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10765 = req_wline & 8'ha8 == req_wset | _GEN_10247; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10766 = req_wline & 8'ha9 == req_wset | _GEN_10248; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10767 = req_wline & 8'haa == req_wset | _GEN_10249; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10768 = req_wline & 8'hab == req_wset | _GEN_10250; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10769 = req_wline & 8'hac == req_wset | _GEN_10251; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10770 = req_wline & 8'had == req_wset | _GEN_10252; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10771 = req_wline & 8'hae == req_wset | _GEN_10253; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10772 = req_wline & 8'haf == req_wset | _GEN_10254; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10773 = req_wline & 8'hb0 == req_wset | _GEN_10255; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10774 = req_wline & 8'hb1 == req_wset | _GEN_10256; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10775 = req_wline & 8'hb2 == req_wset | _GEN_10257; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10776 = req_wline & 8'hb3 == req_wset | _GEN_10258; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10777 = req_wline & 8'hb4 == req_wset | _GEN_10259; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10778 = req_wline & 8'hb5 == req_wset | _GEN_10260; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10779 = req_wline & 8'hb6 == req_wset | _GEN_10261; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10780 = req_wline & 8'hb7 == req_wset | _GEN_10262; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10781 = req_wline & 8'hb8 == req_wset | _GEN_10263; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10782 = req_wline & 8'hb9 == req_wset | _GEN_10264; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10783 = req_wline & 8'hba == req_wset | _GEN_10265; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10784 = req_wline & 8'hbb == req_wset | _GEN_10266; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10785 = req_wline & 8'hbc == req_wset | _GEN_10267; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10786 = req_wline & 8'hbd == req_wset | _GEN_10268; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10787 = req_wline & 8'hbe == req_wset | _GEN_10269; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10788 = req_wline & 8'hbf == req_wset | _GEN_10270; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10789 = req_wline & 8'hc0 == req_wset | _GEN_10271; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10790 = req_wline & 8'hc1 == req_wset | _GEN_10272; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10791 = req_wline & 8'hc2 == req_wset | _GEN_10273; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10792 = req_wline & 8'hc3 == req_wset | _GEN_10274; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10793 = req_wline & 8'hc4 == req_wset | _GEN_10275; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10794 = req_wline & 8'hc5 == req_wset | _GEN_10276; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10795 = req_wline & 8'hc6 == req_wset | _GEN_10277; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10796 = req_wline & 8'hc7 == req_wset | _GEN_10278; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10797 = req_wline & 8'hc8 == req_wset | _GEN_10279; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10798 = req_wline & 8'hc9 == req_wset | _GEN_10280; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10799 = req_wline & 8'hca == req_wset | _GEN_10281; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10800 = req_wline & 8'hcb == req_wset | _GEN_10282; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10801 = req_wline & 8'hcc == req_wset | _GEN_10283; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10802 = req_wline & 8'hcd == req_wset | _GEN_10284; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10803 = req_wline & 8'hce == req_wset | _GEN_10285; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10804 = req_wline & 8'hcf == req_wset | _GEN_10286; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10805 = req_wline & 8'hd0 == req_wset | _GEN_10287; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10806 = req_wline & 8'hd1 == req_wset | _GEN_10288; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10807 = req_wline & 8'hd2 == req_wset | _GEN_10289; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10808 = req_wline & 8'hd3 == req_wset | _GEN_10290; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10809 = req_wline & 8'hd4 == req_wset | _GEN_10291; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10810 = req_wline & 8'hd5 == req_wset | _GEN_10292; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10811 = req_wline & 8'hd6 == req_wset | _GEN_10293; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10812 = req_wline & 8'hd7 == req_wset | _GEN_10294; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10813 = req_wline & 8'hd8 == req_wset | _GEN_10295; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10814 = req_wline & 8'hd9 == req_wset | _GEN_10296; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10815 = req_wline & 8'hda == req_wset | _GEN_10297; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10816 = req_wline & 8'hdb == req_wset | _GEN_10298; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10817 = req_wline & 8'hdc == req_wset | _GEN_10299; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10818 = req_wline & 8'hdd == req_wset | _GEN_10300; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10819 = req_wline & 8'hde == req_wset | _GEN_10301; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10820 = req_wline & 8'hdf == req_wset | _GEN_10302; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10821 = req_wline & 8'he0 == req_wset | _GEN_10303; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10822 = req_wline & 8'he1 == req_wset | _GEN_10304; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10823 = req_wline & 8'he2 == req_wset | _GEN_10305; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10824 = req_wline & 8'he3 == req_wset | _GEN_10306; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10825 = req_wline & 8'he4 == req_wset | _GEN_10307; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10826 = req_wline & 8'he5 == req_wset | _GEN_10308; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10827 = req_wline & 8'he6 == req_wset | _GEN_10309; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10828 = req_wline & 8'he7 == req_wset | _GEN_10310; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10829 = req_wline & 8'he8 == req_wset | _GEN_10311; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10830 = req_wline & 8'he9 == req_wset | _GEN_10312; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10831 = req_wline & 8'hea == req_wset | _GEN_10313; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10832 = req_wline & 8'heb == req_wset | _GEN_10314; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10833 = req_wline & 8'hec == req_wset | _GEN_10315; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10834 = req_wline & 8'hed == req_wset | _GEN_10316; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10835 = req_wline & 8'hee == req_wset | _GEN_10317; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10836 = req_wline & 8'hef == req_wset | _GEN_10318; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10837 = req_wline & 8'hf0 == req_wset | _GEN_10319; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10838 = req_wline & 8'hf1 == req_wset | _GEN_10320; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10839 = req_wline & 8'hf2 == req_wset | _GEN_10321; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10840 = req_wline & 8'hf3 == req_wset | _GEN_10322; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10841 = req_wline & 8'hf4 == req_wset | _GEN_10323; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10842 = req_wline & 8'hf5 == req_wset | _GEN_10324; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10843 = req_wline & 8'hf6 == req_wset | _GEN_10325; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10844 = req_wline & 8'hf7 == req_wset | _GEN_10326; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10845 = req_wline & 8'hf8 == req_wset | _GEN_10327; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10846 = req_wline & 8'hf9 == req_wset | _GEN_10328; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10847 = req_wline & 8'hfa == req_wset | _GEN_10329; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10848 = req_wline & 8'hfb == req_wset | _GEN_10330; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10849 = req_wline & 8'hfc == req_wset | _GEN_10331; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10850 = req_wline & 8'hfd == req_wset | _GEN_10332; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10851 = req_wline & 8'hfe == req_wset | _GEN_10333; // @[dcache.scala 453:{61,61}]
  wire  _GEN_10852 = req_wline & 8'hff == req_wset | _GEN_10334; // @[dcache.scala 453:{61,61}]
  wire  _GEN_17871 = 2'h0 == req_woffset[3:2]; // @[dcache.scala 454:{61,61}]
  wire [7:0] _GEN_10853 = _GEN_16590 & 2'h0 == req_woffset[3:2] ? req_wset : tagv_0_addra; // @[dcache.scala 454:{61,61}]
  wire  _GEN_17873 = 2'h1 == req_woffset[3:2]; // @[dcache.scala 454:{61,61}]
  wire [7:0] _GEN_10854 = _GEN_16590 & 2'h1 == req_woffset[3:2] ? req_wset : tagv_0_addra; // @[dcache.scala 454:{61,61}]
  wire  _GEN_17875 = 2'h2 == req_woffset[3:2]; // @[dcache.scala 454:{61,61}]
  wire [7:0] _GEN_10855 = _GEN_16590 & 2'h2 == req_woffset[3:2] ? req_wset : tagv_0_addra; // @[dcache.scala 454:{61,61}]
  wire  _GEN_17877 = 2'h3 == req_woffset[3:2]; // @[dcache.scala 454:{61,61}]
  wire [7:0] _GEN_10856 = _GEN_16590 & 2'h3 == req_woffset[3:2] ? req_wset : tagv_0_addra; // @[dcache.scala 454:{61,61}]
  wire [7:0] _GEN_10857 = req_wline & 2'h0 == req_woffset[3:2] ? req_wset : tagv_0_addra; // @[dcache.scala 454:{61,61}]
  wire [7:0] _GEN_10858 = req_wline & 2'h1 == req_woffset[3:2] ? req_wset : tagv_0_addra; // @[dcache.scala 454:{61,61}]
  wire [7:0] _GEN_10859 = req_wline & 2'h2 == req_woffset[3:2] ? req_wset : tagv_0_addra; // @[dcache.scala 454:{61,61}]
  wire [7:0] _GEN_10860 = req_wline & 2'h3 == req_woffset[3:2] ? req_wset : tagv_0_addra; // @[dcache.scala 454:{61,61}]
  wire [3:0] _GEN_10861 = _GEN_16590 & _GEN_17871 ? req_wstrb_1 : _GEN_9815; // @[dcache.scala 455:{61,61}]
  wire [3:0] _GEN_10862 = _GEN_16590 & _GEN_17873 ? req_wstrb_1 : _GEN_9816; // @[dcache.scala 455:{61,61}]
  wire [3:0] _GEN_10863 = _GEN_16590 & _GEN_17875 ? req_wstrb_1 : _GEN_9817; // @[dcache.scala 455:{61,61}]
  wire [3:0] _GEN_10864 = _GEN_16590 & _GEN_17877 ? req_wstrb_1 : _GEN_9818; // @[dcache.scala 455:{61,61}]
  wire [3:0] _GEN_10865 = req_wline & _GEN_17871 ? req_wstrb_1 : _GEN_9819; // @[dcache.scala 455:{61,61}]
  wire [3:0] _GEN_10866 = req_wline & _GEN_17873 ? req_wstrb_1 : _GEN_9820; // @[dcache.scala 455:{61,61}]
  wire [3:0] _GEN_10867 = req_wline & _GEN_17875 ? req_wstrb_1 : _GEN_9821; // @[dcache.scala 455:{61,61}]
  wire [3:0] _GEN_10868 = req_wline & _GEN_17877 ? req_wstrb_1 : _GEN_9822; // @[dcache.scala 455:{61,61}]
  wire [31:0] _GEN_10869 = _GEN_16590 & _GEN_17871 ? req_wdata_1 : _GEN_9807; // @[dcache.scala 456:{61,61}]
  wire [31:0] _GEN_10870 = _GEN_16590 & _GEN_17873 ? req_wdata_1 : _GEN_9808; // @[dcache.scala 456:{61,61}]
  wire [31:0] _GEN_10871 = _GEN_16590 & _GEN_17875 ? req_wdata_1 : _GEN_9809; // @[dcache.scala 456:{61,61}]
  wire [31:0] _GEN_10872 = _GEN_16590 & _GEN_17877 ? req_wdata_1 : _GEN_9810; // @[dcache.scala 456:{61,61}]
  wire [31:0] _GEN_10873 = req_wline & _GEN_17871 ? req_wdata_1 : _GEN_9811; // @[dcache.scala 456:{61,61}]
  wire [31:0] _GEN_10874 = req_wline & _GEN_17873 ? req_wdata_1 : _GEN_9812; // @[dcache.scala 456:{61,61}]
  wire [31:0] _GEN_10875 = req_wline & _GEN_17875 ? req_wdata_1 : _GEN_9813; // @[dcache.scala 456:{61,61}]
  wire [31:0] _GEN_10876 = req_wline & _GEN_17877 ? req_wdata_1 : _GEN_9814; // @[dcache.scala 456:{61,61}]
  wire [1:0] _GEN_10878 = _T_53 ? 2'h1 : 2'h0; // @[dcache.scala 469:29 470:31 471:29]
  wire [7:0] _GEN_11392 = 2'h1 == wstate ? _GEN_10853 : tagv_0_addra; // @[dcache.scala 446:19]
  wire [7:0] _GEN_11393 = 2'h1 == wstate ? _GEN_10854 : tagv_0_addra; // @[dcache.scala 446:19]
  wire [7:0] _GEN_11394 = 2'h1 == wstate ? _GEN_10855 : tagv_0_addra; // @[dcache.scala 446:19]
  wire [7:0] _GEN_11395 = 2'h1 == wstate ? _GEN_10856 : tagv_0_addra; // @[dcache.scala 446:19]
  wire [7:0] _GEN_11396 = 2'h1 == wstate ? _GEN_10857 : tagv_0_addra; // @[dcache.scala 446:19]
  wire [7:0] _GEN_11397 = 2'h1 == wstate ? _GEN_10858 : tagv_0_addra; // @[dcache.scala 446:19]
  wire [7:0] _GEN_11398 = 2'h1 == wstate ? _GEN_10859 : tagv_0_addra; // @[dcache.scala 446:19]
  wire [7:0] _GEN_11399 = 2'h1 == wstate ? _GEN_10860 : tagv_0_addra; // @[dcache.scala 446:19]
  wire [3:0] _GEN_11400 = 2'h1 == wstate ? _GEN_10861 : _GEN_9815; // @[dcache.scala 446:19]
  wire [3:0] _GEN_11401 = 2'h1 == wstate ? _GEN_10862 : _GEN_9816; // @[dcache.scala 446:19]
  wire [3:0] _GEN_11402 = 2'h1 == wstate ? _GEN_10863 : _GEN_9817; // @[dcache.scala 446:19]
  wire [3:0] _GEN_11403 = 2'h1 == wstate ? _GEN_10864 : _GEN_9818; // @[dcache.scala 446:19]
  wire [3:0] _GEN_11404 = 2'h1 == wstate ? _GEN_10865 : _GEN_9819; // @[dcache.scala 446:19]
  wire [3:0] _GEN_11405 = 2'h1 == wstate ? _GEN_10866 : _GEN_9820; // @[dcache.scala 446:19]
  wire [3:0] _GEN_11406 = 2'h1 == wstate ? _GEN_10867 : _GEN_9821; // @[dcache.scala 446:19]
  wire [3:0] _GEN_11407 = 2'h1 == wstate ? _GEN_10868 : _GEN_9822; // @[dcache.scala 446:19]
  wire [31:0] _GEN_11408 = 2'h1 == wstate ? _GEN_10869 : _GEN_9807; // @[dcache.scala 446:19]
  wire [31:0] _GEN_11409 = 2'h1 == wstate ? _GEN_10870 : _GEN_9808; // @[dcache.scala 446:19]
  wire [31:0] _GEN_11410 = 2'h1 == wstate ? _GEN_10871 : _GEN_9809; // @[dcache.scala 446:19]
  wire [31:0] _GEN_11411 = 2'h1 == wstate ? _GEN_10872 : _GEN_9810; // @[dcache.scala 446:19]
  wire [31:0] _GEN_11412 = 2'h1 == wstate ? _GEN_10873 : _GEN_9811; // @[dcache.scala 446:19]
  wire [31:0] _GEN_11413 = 2'h1 == wstate ? _GEN_10874 : _GEN_9812; // @[dcache.scala 446:19]
  wire [31:0] _GEN_11414 = 2'h1 == wstate ? _GEN_10875 : _GEN_9813; // @[dcache.scala 446:19]
  wire [31:0] _GEN_11415 = 2'h1 == wstate ? _GEN_10876 : _GEN_9814; // @[dcache.scala 446:19]
  tagv_ram tagv_ram ( // @[dcache.scala 110:49]
    .addra(tagv_ram_addra),
    .clka(tagv_ram_clka),
    .dina(tagv_ram_dina),
    .douta(tagv_ram_douta),
    .wea(tagv_ram_wea)
  );
 tagv_ram tagv_ram_1 ( // @[dcache.scala 110:49]
    .addra(tagv_ram_1_addra),
    .clka(tagv_ram_1_clka),
    .dina(tagv_ram_1_dina),
    .douta(tagv_ram_1_douta),
    .wea(tagv_ram_1_wea)
  );
  data_ram data_ram ( // @[dcache.scala 111:65]
    .addra(data_ram_addra),
    .clka(data_ram_clka),
    .dina(data_ram_dina),
    .douta(data_ram_douta),
    .wea(data_ram_wea)
  );
  data_ram data_ram_1 ( // @[dcache.scala 111:65]
    .addra(data_ram_1_addra),
    .clka(data_ram_1_clka),
    .dina(data_ram_1_dina),
    .douta(data_ram_1_douta),
    .wea(data_ram_1_wea)
  );
  data_ram data_ram_2 ( // @[dcache.scala 111:65]
    .addra(data_ram_2_addra),
    .clka(data_ram_2_clka),
    .dina(data_ram_2_dina),
    .douta(data_ram_2_douta),
    .wea(data_ram_2_wea)
  );
  data_ram data_ram_3 ( // @[dcache.scala 111:65]
    .addra(data_ram_3_addra),
    .clka(data_ram_3_clka),
    .dina(data_ram_3_dina),
    .douta(data_ram_3_douta),
    .wea(data_ram_3_wea)
  );
  data_ram data_ram_4 ( // @[dcache.scala 111:65]
    .addra(data_ram_4_addra),
    .clka(data_ram_4_clka),
    .dina(data_ram_4_dina),
    .douta(data_ram_4_douta),
    .wea(data_ram_4_wea)
  );
  data_ram data_ram_5 ( // @[dcache.scala 111:65]
    .addra(data_ram_5_addra),
    .clka(data_ram_5_clka),
    .dina(data_ram_5_dina),
    .douta(data_ram_5_douta),
    .wea(data_ram_5_wea)
  );
  data_ram data_ram_6 ( // @[dcache.scala 111:65]
    .addra(data_ram_6_addra),
    .clka(data_ram_6_clka),
    .dina(data_ram_6_dina),
    .douta(data_ram_6_douta),
    .wea(data_ram_6_wea)
  );
  data_ram data_ram_7 ( // @[dcache.scala 111:65]
    .addra(data_ram_7_addra),
    .clka(data_ram_7_clka),
    .dina(data_ram_7_dina),
    .douta(data_ram_7_douta),
    .wea(data_ram_7_wea)
  );
  MaxPeriodFibonacciLFSR LFSR_result_prng ( // @[PRNG.scala 91:22]
    .clock(LFSR_result_prng_clock),
    .reset(LFSR_result_prng_reset),
    .io_out_0(LFSR_result_prng_io_out_0),
    .io_out_1(LFSR_result_prng_io_out_1),
    .io_out_2(LFSR_result_prng_io_out_2),
    .io_out_3(LFSR_result_prng_io_out_3),
    .io_out_4(LFSR_result_prng_io_out_4),
    .io_out_5(LFSR_result_prng_io_out_5),
    .io_out_6(LFSR_result_prng_io_out_6),
    .io_out_7(LFSR_result_prng_io_out_7),
    .io_out_8(LFSR_result_prng_io_out_8),
    .io_out_9(LFSR_result_prng_io_out_9),
    .io_out_10(LFSR_result_prng_io_out_10),
    .io_out_11(LFSR_result_prng_io_out_11),
    .io_out_12(LFSR_result_prng_io_out_12),
    .io_out_13(LFSR_result_prng_io_out_13),
    .io_out_14(LFSR_result_prng_io_out_14),
    .io_out_15(LFSR_result_prng_io_out_15)
  );
  assign addr_ok = 3'h0 == state ? _GEN_22 : _GEN_9212; // @[dcache.scala 183:18]
  assign data_ok = 3'h0 == state ? 1'h0 : _GEN_9201; // @[dcache.scala 183:18 157:25]
  assign rdata = 3'h0 == state ? 32'h7777 : _GEN_9193; // @[dcache.scala 183:18 155:25]
  assign rd_req = 3'h0 == state ? 1'h0 : _GEN_9229; // @[dcache.scala 183:18 158:25]
  assign rd_type = 3'h0 == state ? 3'h0 : _GEN_9230; // @[dcache.scala 183:18 159:25]
  assign rd_addr = 3'h0 == state ? 32'h0 : _GEN_9231; // @[dcache.scala 183:18 160:25]
  assign wr_req = 3'h0 == state ? 1'h0 : _GEN_9224; // @[dcache.scala 183:18 161:25]
  assign wr_type = 3'h0 == state ? 3'h0 : _GEN_9227; // @[dcache.scala 183:18 162:25]
  assign wr_addr = 3'h0 == state ? 32'h0 : _GEN_9225; // @[dcache.scala 183:18 163:25]
  assign wr_wstrb = 3'h0 == state ? 4'h0 : _GEN_9228; // @[dcache.scala 183:18 164:25]
  assign wr_data = 3'h0 == state ? 128'h0 : _GEN_9226; // @[dcache.scala 183:18 165:25]
  assign tag_output = 3'h0 == state ? 22'h0 : _GEN_9765; // @[dcache.scala 183:18 98:21]
  assign cache_op_done = 3'h0 == state ? 1'h0 : _GEN_9205; // @[dcache.scala 183:18 97:21]
  assign hit = 3'h0 == state ? 1'h0 : 3'h1 == state & _GEN_72; // @[dcache.scala 183:18 154:25]
  assign tagv_ram_addra = 3'h0 == state ? _GEN_15 : _GEN_9218; // @[dcache.scala 183:18]
  assign tagv_ram_clka = clock; // @[dcache.scala 110:42 142:25]
  assign tagv_ram_dina = 3'h0 == state ? 21'h0 : _GEN_9763; // @[dcache.scala 183:18 143:25]
  assign tagv_ram_wea = 3'h0 == state ? 1'h0 : _GEN_9761; // @[dcache.scala 183:18 144:25]
  assign tagv_ram_1_addra = 3'h0 == state ? _GEN_15 : _GEN_9218; // @[dcache.scala 183:18]
  assign tagv_ram_1_clka = clock; // @[dcache.scala 110:42 142:25]
  assign tagv_ram_1_dina = 3'h0 == state ? 21'h0 : _GEN_9764; // @[dcache.scala 183:18 143:25]
  assign tagv_ram_1_wea = 3'h0 == state ? 1'h0 : _GEN_9762; // @[dcache.scala 183:18 144:25]
  assign data_ram_addra = 2'h0 == wstate ? tagv_0_addra : _GEN_11392; // @[dcache.scala 446:19]
  assign data_ram_clka = clock; // @[dcache.scala 111:58 148:33]
  assign data_ram_dina = 2'h0 == wstate ? _GEN_9807 : _GEN_11408; // @[dcache.scala 446:19]
  assign data_ram_wea = 2'h0 == wstate ? _GEN_9815 : _GEN_11400; // @[dcache.scala 446:19]
  assign data_ram_1_addra = 2'h0 == wstate ? tagv_0_addra : _GEN_11393; // @[dcache.scala 446:19]
  assign data_ram_1_clka = clock; // @[dcache.scala 111:58 148:33]
  assign data_ram_1_dina = 2'h0 == wstate ? _GEN_9808 : _GEN_11409; // @[dcache.scala 446:19]
  assign data_ram_1_wea = 2'h0 == wstate ? _GEN_9816 : _GEN_11401; // @[dcache.scala 446:19]
  assign data_ram_2_addra = 2'h0 == wstate ? tagv_0_addra : _GEN_11394; // @[dcache.scala 446:19]
  assign data_ram_2_clka = clock; // @[dcache.scala 111:58 148:33]
  assign data_ram_2_dina = 2'h0 == wstate ? _GEN_9809 : _GEN_11410; // @[dcache.scala 446:19]
  assign data_ram_2_wea = 2'h0 == wstate ? _GEN_9817 : _GEN_11402; // @[dcache.scala 446:19]
  assign data_ram_3_addra = 2'h0 == wstate ? tagv_0_addra : _GEN_11395; // @[dcache.scala 446:19]
  assign data_ram_3_clka = clock; // @[dcache.scala 111:58 148:33]
  assign data_ram_3_dina = 2'h0 == wstate ? _GEN_9810 : _GEN_11411; // @[dcache.scala 446:19]
  assign data_ram_3_wea = 2'h0 == wstate ? _GEN_9818 : _GEN_11403; // @[dcache.scala 446:19]
  assign data_ram_4_addra = 2'h0 == wstate ? tagv_0_addra : _GEN_11396; // @[dcache.scala 446:19]
  assign data_ram_4_clka = clock; // @[dcache.scala 111:58 148:33]
  assign data_ram_4_dina = 2'h0 == wstate ? _GEN_9811 : _GEN_11412; // @[dcache.scala 446:19]
  assign data_ram_4_wea = 2'h0 == wstate ? _GEN_9819 : _GEN_11404; // @[dcache.scala 446:19]
  assign data_ram_5_addra = 2'h0 == wstate ? tagv_0_addra : _GEN_11397; // @[dcache.scala 446:19]
  assign data_ram_5_clka = clock; // @[dcache.scala 111:58 148:33]
  assign data_ram_5_dina = 2'h0 == wstate ? _GEN_9812 : _GEN_11413; // @[dcache.scala 446:19]
  assign data_ram_5_wea = 2'h0 == wstate ? _GEN_9820 : _GEN_11405; // @[dcache.scala 446:19]
  assign data_ram_6_addra = 2'h0 == wstate ? tagv_0_addra : _GEN_11398; // @[dcache.scala 446:19]
  assign data_ram_6_clka = clock; // @[dcache.scala 111:58 148:33]
  assign data_ram_6_dina = 2'h0 == wstate ? _GEN_9813 : _GEN_11414; // @[dcache.scala 446:19]
  assign data_ram_6_wea = 2'h0 == wstate ? _GEN_9821 : _GEN_11406; // @[dcache.scala 446:19]
  assign data_ram_7_addra = 2'h0 == wstate ? tagv_0_addra : _GEN_11399; // @[dcache.scala 446:19]
  assign data_ram_7_clka = clock; // @[dcache.scala 111:58 148:33]
  assign data_ram_7_dina = 2'h0 == wstate ? _GEN_9814 : _GEN_11415; // @[dcache.scala 446:19]
  assign data_ram_7_wea = 2'h0 == wstate ? _GEN_9822 : _GEN_11407; // @[dcache.scala 446:19]
  assign LFSR_result_prng_clock = clock;
  assign LFSR_result_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[dcache.scala 89:38]
      cacheInst_r <= 1'h0; // @[dcache.scala 89:38]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        cacheInst_r <= cache_op_en; // @[dcache.scala 191:33]
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (cacheInst_r) begin // @[dcache.scala 255:30]
        cacheInst_r <= _GEN_93;
      end
    end else if (!(3'h2 == state)) begin // @[dcache.scala 183:18]
      cacheInst_r <= _GEN_8629;
    end
    if (reset) begin // @[dcache.scala 90:38]
      invalidate <= 1'h0; // @[dcache.scala 90:38]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        invalidate <= cacheOperation_0; // @[dcache.scala 192:33]
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (cacheInst_r) begin // @[dcache.scala 255:30]
        invalidate <= _GEN_94;
      end
    end else if (!(3'h2 == state)) begin // @[dcache.scala 183:18]
      invalidate <= _GEN_8630;
    end
    if (reset) begin // @[dcache.scala 91:38]
      loadTag <= 1'h0; // @[dcache.scala 91:38]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        if (_cacheOperation_T_1) begin // @[Lookup.scala 34:39]
          loadTag <= 1'h0;
        end else begin
          loadTag <= _cacheOperation_T_3;
        end
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (cacheInst_r) begin // @[dcache.scala 255:30]
        loadTag <= _GEN_98;
      end
    end else if (!(3'h2 == state)) begin // @[dcache.scala 183:18]
      loadTag <= _GEN_8634;
    end
    if (reset) begin // @[dcache.scala 92:38]
      storeTag <= 1'h0; // @[dcache.scala 92:38]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        if (_cacheOperation_T_1) begin // @[Lookup.scala 34:39]
          storeTag <= 1'h0;
        end else begin
          storeTag <= _cacheOperation_T_36;
        end
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (cacheInst_r) begin // @[dcache.scala 255:30]
        storeTag <= _GEN_97;
      end
    end else if (!(3'h2 == state)) begin // @[dcache.scala 183:18]
      storeTag <= _GEN_8633;
    end
    if (reset) begin // @[dcache.scala 93:38]
      writeBack <= 1'h0; // @[dcache.scala 93:38]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        writeBack <= cacheOperation_3; // @[dcache.scala 195:33]
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (cacheInst_r) begin // @[dcache.scala 255:30]
        writeBack <= _GEN_96;
      end
    end else if (!(3'h2 == state)) begin // @[dcache.scala 183:18]
      writeBack <= _GEN_8632;
    end
    if (reset) begin // @[dcache.scala 94:38]
      indexOnly <= 1'h0; // @[dcache.scala 94:38]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        indexOnly <= cacheOperation_4; // @[dcache.scala 196:33]
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (cacheInst_r) begin // @[dcache.scala 255:30]
        indexOnly <= _GEN_95;
      end
    end else if (!(3'h2 == state)) begin // @[dcache.scala 183:18]
      indexOnly <= _GEN_8631;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_0 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_0 <= _GEN_9823;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_0 <= _GEN_10341;
    end else begin
      dirty_0_0 <= _GEN_9823;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_1 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_1 <= _GEN_9824;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_1 <= _GEN_10342;
    end else begin
      dirty_0_1 <= _GEN_9824;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_2 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_2 <= _GEN_9825;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_2 <= _GEN_10343;
    end else begin
      dirty_0_2 <= _GEN_9825;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_3 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_3 <= _GEN_9826;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_3 <= _GEN_10344;
    end else begin
      dirty_0_3 <= _GEN_9826;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_4 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_4 <= _GEN_9827;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_4 <= _GEN_10345;
    end else begin
      dirty_0_4 <= _GEN_9827;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_5 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_5 <= _GEN_9828;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_5 <= _GEN_10346;
    end else begin
      dirty_0_5 <= _GEN_9828;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_6 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_6 <= _GEN_9829;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_6 <= _GEN_10347;
    end else begin
      dirty_0_6 <= _GEN_9829;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_7 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_7 <= _GEN_9830;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_7 <= _GEN_10348;
    end else begin
      dirty_0_7 <= _GEN_9830;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_8 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_8 <= _GEN_9831;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_8 <= _GEN_10349;
    end else begin
      dirty_0_8 <= _GEN_9831;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_9 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_9 <= _GEN_9832;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_9 <= _GEN_10350;
    end else begin
      dirty_0_9 <= _GEN_9832;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_10 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_10 <= _GEN_9833;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_10 <= _GEN_10351;
    end else begin
      dirty_0_10 <= _GEN_9833;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_11 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_11 <= _GEN_9834;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_11 <= _GEN_10352;
    end else begin
      dirty_0_11 <= _GEN_9834;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_12 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_12 <= _GEN_9835;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_12 <= _GEN_10353;
    end else begin
      dirty_0_12 <= _GEN_9835;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_13 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_13 <= _GEN_9836;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_13 <= _GEN_10354;
    end else begin
      dirty_0_13 <= _GEN_9836;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_14 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_14 <= _GEN_9837;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_14 <= _GEN_10355;
    end else begin
      dirty_0_14 <= _GEN_9837;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_15 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_15 <= _GEN_9838;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_15 <= _GEN_10356;
    end else begin
      dirty_0_15 <= _GEN_9838;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_16 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_16 <= _GEN_9839;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_16 <= _GEN_10357;
    end else begin
      dirty_0_16 <= _GEN_9839;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_17 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_17 <= _GEN_9840;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_17 <= _GEN_10358;
    end else begin
      dirty_0_17 <= _GEN_9840;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_18 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_18 <= _GEN_9841;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_18 <= _GEN_10359;
    end else begin
      dirty_0_18 <= _GEN_9841;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_19 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_19 <= _GEN_9842;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_19 <= _GEN_10360;
    end else begin
      dirty_0_19 <= _GEN_9842;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_20 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_20 <= _GEN_9843;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_20 <= _GEN_10361;
    end else begin
      dirty_0_20 <= _GEN_9843;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_21 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_21 <= _GEN_9844;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_21 <= _GEN_10362;
    end else begin
      dirty_0_21 <= _GEN_9844;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_22 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_22 <= _GEN_9845;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_22 <= _GEN_10363;
    end else begin
      dirty_0_22 <= _GEN_9845;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_23 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_23 <= _GEN_9846;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_23 <= _GEN_10364;
    end else begin
      dirty_0_23 <= _GEN_9846;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_24 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_24 <= _GEN_9847;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_24 <= _GEN_10365;
    end else begin
      dirty_0_24 <= _GEN_9847;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_25 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_25 <= _GEN_9848;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_25 <= _GEN_10366;
    end else begin
      dirty_0_25 <= _GEN_9848;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_26 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_26 <= _GEN_9849;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_26 <= _GEN_10367;
    end else begin
      dirty_0_26 <= _GEN_9849;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_27 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_27 <= _GEN_9850;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_27 <= _GEN_10368;
    end else begin
      dirty_0_27 <= _GEN_9850;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_28 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_28 <= _GEN_9851;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_28 <= _GEN_10369;
    end else begin
      dirty_0_28 <= _GEN_9851;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_29 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_29 <= _GEN_9852;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_29 <= _GEN_10370;
    end else begin
      dirty_0_29 <= _GEN_9852;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_30 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_30 <= _GEN_9853;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_30 <= _GEN_10371;
    end else begin
      dirty_0_30 <= _GEN_9853;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_31 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_31 <= _GEN_9854;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_31 <= _GEN_10372;
    end else begin
      dirty_0_31 <= _GEN_9854;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_32 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_32 <= _GEN_9855;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_32 <= _GEN_10373;
    end else begin
      dirty_0_32 <= _GEN_9855;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_33 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_33 <= _GEN_9856;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_33 <= _GEN_10374;
    end else begin
      dirty_0_33 <= _GEN_9856;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_34 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_34 <= _GEN_9857;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_34 <= _GEN_10375;
    end else begin
      dirty_0_34 <= _GEN_9857;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_35 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_35 <= _GEN_9858;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_35 <= _GEN_10376;
    end else begin
      dirty_0_35 <= _GEN_9858;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_36 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_36 <= _GEN_9859;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_36 <= _GEN_10377;
    end else begin
      dirty_0_36 <= _GEN_9859;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_37 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_37 <= _GEN_9860;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_37 <= _GEN_10378;
    end else begin
      dirty_0_37 <= _GEN_9860;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_38 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_38 <= _GEN_9861;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_38 <= _GEN_10379;
    end else begin
      dirty_0_38 <= _GEN_9861;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_39 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_39 <= _GEN_9862;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_39 <= _GEN_10380;
    end else begin
      dirty_0_39 <= _GEN_9862;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_40 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_40 <= _GEN_9863;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_40 <= _GEN_10381;
    end else begin
      dirty_0_40 <= _GEN_9863;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_41 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_41 <= _GEN_9864;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_41 <= _GEN_10382;
    end else begin
      dirty_0_41 <= _GEN_9864;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_42 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_42 <= _GEN_9865;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_42 <= _GEN_10383;
    end else begin
      dirty_0_42 <= _GEN_9865;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_43 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_43 <= _GEN_9866;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_43 <= _GEN_10384;
    end else begin
      dirty_0_43 <= _GEN_9866;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_44 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_44 <= _GEN_9867;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_44 <= _GEN_10385;
    end else begin
      dirty_0_44 <= _GEN_9867;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_45 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_45 <= _GEN_9868;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_45 <= _GEN_10386;
    end else begin
      dirty_0_45 <= _GEN_9868;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_46 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_46 <= _GEN_9869;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_46 <= _GEN_10387;
    end else begin
      dirty_0_46 <= _GEN_9869;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_47 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_47 <= _GEN_9870;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_47 <= _GEN_10388;
    end else begin
      dirty_0_47 <= _GEN_9870;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_48 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_48 <= _GEN_9871;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_48 <= _GEN_10389;
    end else begin
      dirty_0_48 <= _GEN_9871;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_49 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_49 <= _GEN_9872;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_49 <= _GEN_10390;
    end else begin
      dirty_0_49 <= _GEN_9872;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_50 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_50 <= _GEN_9873;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_50 <= _GEN_10391;
    end else begin
      dirty_0_50 <= _GEN_9873;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_51 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_51 <= _GEN_9874;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_51 <= _GEN_10392;
    end else begin
      dirty_0_51 <= _GEN_9874;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_52 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_52 <= _GEN_9875;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_52 <= _GEN_10393;
    end else begin
      dirty_0_52 <= _GEN_9875;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_53 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_53 <= _GEN_9876;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_53 <= _GEN_10394;
    end else begin
      dirty_0_53 <= _GEN_9876;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_54 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_54 <= _GEN_9877;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_54 <= _GEN_10395;
    end else begin
      dirty_0_54 <= _GEN_9877;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_55 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_55 <= _GEN_9878;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_55 <= _GEN_10396;
    end else begin
      dirty_0_55 <= _GEN_9878;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_56 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_56 <= _GEN_9879;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_56 <= _GEN_10397;
    end else begin
      dirty_0_56 <= _GEN_9879;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_57 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_57 <= _GEN_9880;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_57 <= _GEN_10398;
    end else begin
      dirty_0_57 <= _GEN_9880;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_58 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_58 <= _GEN_9881;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_58 <= _GEN_10399;
    end else begin
      dirty_0_58 <= _GEN_9881;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_59 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_59 <= _GEN_9882;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_59 <= _GEN_10400;
    end else begin
      dirty_0_59 <= _GEN_9882;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_60 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_60 <= _GEN_9883;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_60 <= _GEN_10401;
    end else begin
      dirty_0_60 <= _GEN_9883;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_61 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_61 <= _GEN_9884;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_61 <= _GEN_10402;
    end else begin
      dirty_0_61 <= _GEN_9884;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_62 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_62 <= _GEN_9885;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_62 <= _GEN_10403;
    end else begin
      dirty_0_62 <= _GEN_9885;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_63 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_63 <= _GEN_9886;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_63 <= _GEN_10404;
    end else begin
      dirty_0_63 <= _GEN_9886;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_64 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_64 <= _GEN_9887;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_64 <= _GEN_10405;
    end else begin
      dirty_0_64 <= _GEN_9887;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_65 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_65 <= _GEN_9888;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_65 <= _GEN_10406;
    end else begin
      dirty_0_65 <= _GEN_9888;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_66 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_66 <= _GEN_9889;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_66 <= _GEN_10407;
    end else begin
      dirty_0_66 <= _GEN_9889;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_67 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_67 <= _GEN_9890;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_67 <= _GEN_10408;
    end else begin
      dirty_0_67 <= _GEN_9890;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_68 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_68 <= _GEN_9891;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_68 <= _GEN_10409;
    end else begin
      dirty_0_68 <= _GEN_9891;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_69 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_69 <= _GEN_9892;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_69 <= _GEN_10410;
    end else begin
      dirty_0_69 <= _GEN_9892;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_70 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_70 <= _GEN_9893;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_70 <= _GEN_10411;
    end else begin
      dirty_0_70 <= _GEN_9893;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_71 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_71 <= _GEN_9894;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_71 <= _GEN_10412;
    end else begin
      dirty_0_71 <= _GEN_9894;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_72 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_72 <= _GEN_9895;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_72 <= _GEN_10413;
    end else begin
      dirty_0_72 <= _GEN_9895;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_73 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_73 <= _GEN_9896;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_73 <= _GEN_10414;
    end else begin
      dirty_0_73 <= _GEN_9896;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_74 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_74 <= _GEN_9897;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_74 <= _GEN_10415;
    end else begin
      dirty_0_74 <= _GEN_9897;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_75 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_75 <= _GEN_9898;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_75 <= _GEN_10416;
    end else begin
      dirty_0_75 <= _GEN_9898;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_76 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_76 <= _GEN_9899;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_76 <= _GEN_10417;
    end else begin
      dirty_0_76 <= _GEN_9899;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_77 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_77 <= _GEN_9900;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_77 <= _GEN_10418;
    end else begin
      dirty_0_77 <= _GEN_9900;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_78 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_78 <= _GEN_9901;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_78 <= _GEN_10419;
    end else begin
      dirty_0_78 <= _GEN_9901;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_79 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_79 <= _GEN_9902;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_79 <= _GEN_10420;
    end else begin
      dirty_0_79 <= _GEN_9902;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_80 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_80 <= _GEN_9903;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_80 <= _GEN_10421;
    end else begin
      dirty_0_80 <= _GEN_9903;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_81 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_81 <= _GEN_9904;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_81 <= _GEN_10422;
    end else begin
      dirty_0_81 <= _GEN_9904;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_82 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_82 <= _GEN_9905;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_82 <= _GEN_10423;
    end else begin
      dirty_0_82 <= _GEN_9905;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_83 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_83 <= _GEN_9906;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_83 <= _GEN_10424;
    end else begin
      dirty_0_83 <= _GEN_9906;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_84 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_84 <= _GEN_9907;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_84 <= _GEN_10425;
    end else begin
      dirty_0_84 <= _GEN_9907;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_85 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_85 <= _GEN_9908;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_85 <= _GEN_10426;
    end else begin
      dirty_0_85 <= _GEN_9908;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_86 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_86 <= _GEN_9909;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_86 <= _GEN_10427;
    end else begin
      dirty_0_86 <= _GEN_9909;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_87 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_87 <= _GEN_9910;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_87 <= _GEN_10428;
    end else begin
      dirty_0_87 <= _GEN_9910;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_88 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_88 <= _GEN_9911;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_88 <= _GEN_10429;
    end else begin
      dirty_0_88 <= _GEN_9911;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_89 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_89 <= _GEN_9912;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_89 <= _GEN_10430;
    end else begin
      dirty_0_89 <= _GEN_9912;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_90 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_90 <= _GEN_9913;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_90 <= _GEN_10431;
    end else begin
      dirty_0_90 <= _GEN_9913;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_91 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_91 <= _GEN_9914;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_91 <= _GEN_10432;
    end else begin
      dirty_0_91 <= _GEN_9914;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_92 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_92 <= _GEN_9915;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_92 <= _GEN_10433;
    end else begin
      dirty_0_92 <= _GEN_9915;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_93 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_93 <= _GEN_9916;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_93 <= _GEN_10434;
    end else begin
      dirty_0_93 <= _GEN_9916;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_94 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_94 <= _GEN_9917;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_94 <= _GEN_10435;
    end else begin
      dirty_0_94 <= _GEN_9917;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_95 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_95 <= _GEN_9918;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_95 <= _GEN_10436;
    end else begin
      dirty_0_95 <= _GEN_9918;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_96 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_96 <= _GEN_9919;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_96 <= _GEN_10437;
    end else begin
      dirty_0_96 <= _GEN_9919;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_97 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_97 <= _GEN_9920;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_97 <= _GEN_10438;
    end else begin
      dirty_0_97 <= _GEN_9920;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_98 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_98 <= _GEN_9921;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_98 <= _GEN_10439;
    end else begin
      dirty_0_98 <= _GEN_9921;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_99 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_99 <= _GEN_9922;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_99 <= _GEN_10440;
    end else begin
      dirty_0_99 <= _GEN_9922;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_100 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_100 <= _GEN_9923;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_100 <= _GEN_10441;
    end else begin
      dirty_0_100 <= _GEN_9923;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_101 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_101 <= _GEN_9924;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_101 <= _GEN_10442;
    end else begin
      dirty_0_101 <= _GEN_9924;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_102 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_102 <= _GEN_9925;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_102 <= _GEN_10443;
    end else begin
      dirty_0_102 <= _GEN_9925;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_103 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_103 <= _GEN_9926;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_103 <= _GEN_10444;
    end else begin
      dirty_0_103 <= _GEN_9926;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_104 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_104 <= _GEN_9927;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_104 <= _GEN_10445;
    end else begin
      dirty_0_104 <= _GEN_9927;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_105 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_105 <= _GEN_9928;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_105 <= _GEN_10446;
    end else begin
      dirty_0_105 <= _GEN_9928;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_106 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_106 <= _GEN_9929;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_106 <= _GEN_10447;
    end else begin
      dirty_0_106 <= _GEN_9929;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_107 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_107 <= _GEN_9930;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_107 <= _GEN_10448;
    end else begin
      dirty_0_107 <= _GEN_9930;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_108 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_108 <= _GEN_9931;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_108 <= _GEN_10449;
    end else begin
      dirty_0_108 <= _GEN_9931;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_109 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_109 <= _GEN_9932;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_109 <= _GEN_10450;
    end else begin
      dirty_0_109 <= _GEN_9932;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_110 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_110 <= _GEN_9933;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_110 <= _GEN_10451;
    end else begin
      dirty_0_110 <= _GEN_9933;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_111 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_111 <= _GEN_9934;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_111 <= _GEN_10452;
    end else begin
      dirty_0_111 <= _GEN_9934;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_112 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_112 <= _GEN_9935;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_112 <= _GEN_10453;
    end else begin
      dirty_0_112 <= _GEN_9935;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_113 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_113 <= _GEN_9936;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_113 <= _GEN_10454;
    end else begin
      dirty_0_113 <= _GEN_9936;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_114 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_114 <= _GEN_9937;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_114 <= _GEN_10455;
    end else begin
      dirty_0_114 <= _GEN_9937;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_115 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_115 <= _GEN_9938;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_115 <= _GEN_10456;
    end else begin
      dirty_0_115 <= _GEN_9938;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_116 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_116 <= _GEN_9939;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_116 <= _GEN_10457;
    end else begin
      dirty_0_116 <= _GEN_9939;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_117 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_117 <= _GEN_9940;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_117 <= _GEN_10458;
    end else begin
      dirty_0_117 <= _GEN_9940;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_118 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_118 <= _GEN_9941;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_118 <= _GEN_10459;
    end else begin
      dirty_0_118 <= _GEN_9941;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_119 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_119 <= _GEN_9942;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_119 <= _GEN_10460;
    end else begin
      dirty_0_119 <= _GEN_9942;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_120 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_120 <= _GEN_9943;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_120 <= _GEN_10461;
    end else begin
      dirty_0_120 <= _GEN_9943;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_121 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_121 <= _GEN_9944;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_121 <= _GEN_10462;
    end else begin
      dirty_0_121 <= _GEN_9944;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_122 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_122 <= _GEN_9945;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_122 <= _GEN_10463;
    end else begin
      dirty_0_122 <= _GEN_9945;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_123 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_123 <= _GEN_9946;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_123 <= _GEN_10464;
    end else begin
      dirty_0_123 <= _GEN_9946;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_124 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_124 <= _GEN_9947;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_124 <= _GEN_10465;
    end else begin
      dirty_0_124 <= _GEN_9947;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_125 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_125 <= _GEN_9948;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_125 <= _GEN_10466;
    end else begin
      dirty_0_125 <= _GEN_9948;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_126 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_126 <= _GEN_9949;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_126 <= _GEN_10467;
    end else begin
      dirty_0_126 <= _GEN_9949;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_127 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_127 <= _GEN_9950;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_127 <= _GEN_10468;
    end else begin
      dirty_0_127 <= _GEN_9950;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_128 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_128 <= _GEN_9951;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_128 <= _GEN_10469;
    end else begin
      dirty_0_128 <= _GEN_9951;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_129 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_129 <= _GEN_9952;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_129 <= _GEN_10470;
    end else begin
      dirty_0_129 <= _GEN_9952;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_130 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_130 <= _GEN_9953;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_130 <= _GEN_10471;
    end else begin
      dirty_0_130 <= _GEN_9953;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_131 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_131 <= _GEN_9954;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_131 <= _GEN_10472;
    end else begin
      dirty_0_131 <= _GEN_9954;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_132 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_132 <= _GEN_9955;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_132 <= _GEN_10473;
    end else begin
      dirty_0_132 <= _GEN_9955;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_133 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_133 <= _GEN_9956;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_133 <= _GEN_10474;
    end else begin
      dirty_0_133 <= _GEN_9956;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_134 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_134 <= _GEN_9957;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_134 <= _GEN_10475;
    end else begin
      dirty_0_134 <= _GEN_9957;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_135 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_135 <= _GEN_9958;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_135 <= _GEN_10476;
    end else begin
      dirty_0_135 <= _GEN_9958;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_136 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_136 <= _GEN_9959;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_136 <= _GEN_10477;
    end else begin
      dirty_0_136 <= _GEN_9959;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_137 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_137 <= _GEN_9960;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_137 <= _GEN_10478;
    end else begin
      dirty_0_137 <= _GEN_9960;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_138 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_138 <= _GEN_9961;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_138 <= _GEN_10479;
    end else begin
      dirty_0_138 <= _GEN_9961;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_139 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_139 <= _GEN_9962;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_139 <= _GEN_10480;
    end else begin
      dirty_0_139 <= _GEN_9962;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_140 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_140 <= _GEN_9963;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_140 <= _GEN_10481;
    end else begin
      dirty_0_140 <= _GEN_9963;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_141 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_141 <= _GEN_9964;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_141 <= _GEN_10482;
    end else begin
      dirty_0_141 <= _GEN_9964;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_142 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_142 <= _GEN_9965;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_142 <= _GEN_10483;
    end else begin
      dirty_0_142 <= _GEN_9965;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_143 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_143 <= _GEN_9966;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_143 <= _GEN_10484;
    end else begin
      dirty_0_143 <= _GEN_9966;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_144 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_144 <= _GEN_9967;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_144 <= _GEN_10485;
    end else begin
      dirty_0_144 <= _GEN_9967;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_145 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_145 <= _GEN_9968;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_145 <= _GEN_10486;
    end else begin
      dirty_0_145 <= _GEN_9968;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_146 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_146 <= _GEN_9969;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_146 <= _GEN_10487;
    end else begin
      dirty_0_146 <= _GEN_9969;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_147 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_147 <= _GEN_9970;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_147 <= _GEN_10488;
    end else begin
      dirty_0_147 <= _GEN_9970;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_148 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_148 <= _GEN_9971;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_148 <= _GEN_10489;
    end else begin
      dirty_0_148 <= _GEN_9971;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_149 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_149 <= _GEN_9972;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_149 <= _GEN_10490;
    end else begin
      dirty_0_149 <= _GEN_9972;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_150 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_150 <= _GEN_9973;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_150 <= _GEN_10491;
    end else begin
      dirty_0_150 <= _GEN_9973;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_151 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_151 <= _GEN_9974;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_151 <= _GEN_10492;
    end else begin
      dirty_0_151 <= _GEN_9974;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_152 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_152 <= _GEN_9975;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_152 <= _GEN_10493;
    end else begin
      dirty_0_152 <= _GEN_9975;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_153 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_153 <= _GEN_9976;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_153 <= _GEN_10494;
    end else begin
      dirty_0_153 <= _GEN_9976;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_154 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_154 <= _GEN_9977;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_154 <= _GEN_10495;
    end else begin
      dirty_0_154 <= _GEN_9977;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_155 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_155 <= _GEN_9978;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_155 <= _GEN_10496;
    end else begin
      dirty_0_155 <= _GEN_9978;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_156 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_156 <= _GEN_9979;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_156 <= _GEN_10497;
    end else begin
      dirty_0_156 <= _GEN_9979;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_157 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_157 <= _GEN_9980;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_157 <= _GEN_10498;
    end else begin
      dirty_0_157 <= _GEN_9980;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_158 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_158 <= _GEN_9981;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_158 <= _GEN_10499;
    end else begin
      dirty_0_158 <= _GEN_9981;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_159 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_159 <= _GEN_9982;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_159 <= _GEN_10500;
    end else begin
      dirty_0_159 <= _GEN_9982;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_160 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_160 <= _GEN_9983;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_160 <= _GEN_10501;
    end else begin
      dirty_0_160 <= _GEN_9983;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_161 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_161 <= _GEN_9984;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_161 <= _GEN_10502;
    end else begin
      dirty_0_161 <= _GEN_9984;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_162 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_162 <= _GEN_9985;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_162 <= _GEN_10503;
    end else begin
      dirty_0_162 <= _GEN_9985;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_163 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_163 <= _GEN_9986;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_163 <= _GEN_10504;
    end else begin
      dirty_0_163 <= _GEN_9986;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_164 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_164 <= _GEN_9987;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_164 <= _GEN_10505;
    end else begin
      dirty_0_164 <= _GEN_9987;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_165 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_165 <= _GEN_9988;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_165 <= _GEN_10506;
    end else begin
      dirty_0_165 <= _GEN_9988;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_166 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_166 <= _GEN_9989;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_166 <= _GEN_10507;
    end else begin
      dirty_0_166 <= _GEN_9989;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_167 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_167 <= _GEN_9990;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_167 <= _GEN_10508;
    end else begin
      dirty_0_167 <= _GEN_9990;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_168 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_168 <= _GEN_9991;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_168 <= _GEN_10509;
    end else begin
      dirty_0_168 <= _GEN_9991;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_169 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_169 <= _GEN_9992;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_169 <= _GEN_10510;
    end else begin
      dirty_0_169 <= _GEN_9992;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_170 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_170 <= _GEN_9993;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_170 <= _GEN_10511;
    end else begin
      dirty_0_170 <= _GEN_9993;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_171 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_171 <= _GEN_9994;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_171 <= _GEN_10512;
    end else begin
      dirty_0_171 <= _GEN_9994;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_172 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_172 <= _GEN_9995;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_172 <= _GEN_10513;
    end else begin
      dirty_0_172 <= _GEN_9995;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_173 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_173 <= _GEN_9996;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_173 <= _GEN_10514;
    end else begin
      dirty_0_173 <= _GEN_9996;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_174 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_174 <= _GEN_9997;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_174 <= _GEN_10515;
    end else begin
      dirty_0_174 <= _GEN_9997;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_175 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_175 <= _GEN_9998;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_175 <= _GEN_10516;
    end else begin
      dirty_0_175 <= _GEN_9998;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_176 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_176 <= _GEN_9999;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_176 <= _GEN_10517;
    end else begin
      dirty_0_176 <= _GEN_9999;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_177 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_177 <= _GEN_10000;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_177 <= _GEN_10518;
    end else begin
      dirty_0_177 <= _GEN_10000;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_178 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_178 <= _GEN_10001;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_178 <= _GEN_10519;
    end else begin
      dirty_0_178 <= _GEN_10001;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_179 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_179 <= _GEN_10002;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_179 <= _GEN_10520;
    end else begin
      dirty_0_179 <= _GEN_10002;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_180 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_180 <= _GEN_10003;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_180 <= _GEN_10521;
    end else begin
      dirty_0_180 <= _GEN_10003;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_181 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_181 <= _GEN_10004;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_181 <= _GEN_10522;
    end else begin
      dirty_0_181 <= _GEN_10004;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_182 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_182 <= _GEN_10005;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_182 <= _GEN_10523;
    end else begin
      dirty_0_182 <= _GEN_10005;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_183 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_183 <= _GEN_10006;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_183 <= _GEN_10524;
    end else begin
      dirty_0_183 <= _GEN_10006;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_184 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_184 <= _GEN_10007;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_184 <= _GEN_10525;
    end else begin
      dirty_0_184 <= _GEN_10007;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_185 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_185 <= _GEN_10008;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_185 <= _GEN_10526;
    end else begin
      dirty_0_185 <= _GEN_10008;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_186 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_186 <= _GEN_10009;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_186 <= _GEN_10527;
    end else begin
      dirty_0_186 <= _GEN_10009;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_187 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_187 <= _GEN_10010;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_187 <= _GEN_10528;
    end else begin
      dirty_0_187 <= _GEN_10010;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_188 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_188 <= _GEN_10011;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_188 <= _GEN_10529;
    end else begin
      dirty_0_188 <= _GEN_10011;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_189 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_189 <= _GEN_10012;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_189 <= _GEN_10530;
    end else begin
      dirty_0_189 <= _GEN_10012;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_190 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_190 <= _GEN_10013;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_190 <= _GEN_10531;
    end else begin
      dirty_0_190 <= _GEN_10013;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_191 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_191 <= _GEN_10014;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_191 <= _GEN_10532;
    end else begin
      dirty_0_191 <= _GEN_10014;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_192 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_192 <= _GEN_10015;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_192 <= _GEN_10533;
    end else begin
      dirty_0_192 <= _GEN_10015;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_193 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_193 <= _GEN_10016;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_193 <= _GEN_10534;
    end else begin
      dirty_0_193 <= _GEN_10016;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_194 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_194 <= _GEN_10017;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_194 <= _GEN_10535;
    end else begin
      dirty_0_194 <= _GEN_10017;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_195 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_195 <= _GEN_10018;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_195 <= _GEN_10536;
    end else begin
      dirty_0_195 <= _GEN_10018;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_196 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_196 <= _GEN_10019;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_196 <= _GEN_10537;
    end else begin
      dirty_0_196 <= _GEN_10019;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_197 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_197 <= _GEN_10020;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_197 <= _GEN_10538;
    end else begin
      dirty_0_197 <= _GEN_10020;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_198 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_198 <= _GEN_10021;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_198 <= _GEN_10539;
    end else begin
      dirty_0_198 <= _GEN_10021;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_199 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_199 <= _GEN_10022;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_199 <= _GEN_10540;
    end else begin
      dirty_0_199 <= _GEN_10022;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_200 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_200 <= _GEN_10023;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_200 <= _GEN_10541;
    end else begin
      dirty_0_200 <= _GEN_10023;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_201 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_201 <= _GEN_10024;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_201 <= _GEN_10542;
    end else begin
      dirty_0_201 <= _GEN_10024;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_202 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_202 <= _GEN_10025;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_202 <= _GEN_10543;
    end else begin
      dirty_0_202 <= _GEN_10025;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_203 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_203 <= _GEN_10026;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_203 <= _GEN_10544;
    end else begin
      dirty_0_203 <= _GEN_10026;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_204 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_204 <= _GEN_10027;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_204 <= _GEN_10545;
    end else begin
      dirty_0_204 <= _GEN_10027;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_205 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_205 <= _GEN_10028;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_205 <= _GEN_10546;
    end else begin
      dirty_0_205 <= _GEN_10028;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_206 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_206 <= _GEN_10029;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_206 <= _GEN_10547;
    end else begin
      dirty_0_206 <= _GEN_10029;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_207 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_207 <= _GEN_10030;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_207 <= _GEN_10548;
    end else begin
      dirty_0_207 <= _GEN_10030;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_208 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_208 <= _GEN_10031;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_208 <= _GEN_10549;
    end else begin
      dirty_0_208 <= _GEN_10031;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_209 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_209 <= _GEN_10032;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_209 <= _GEN_10550;
    end else begin
      dirty_0_209 <= _GEN_10032;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_210 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_210 <= _GEN_10033;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_210 <= _GEN_10551;
    end else begin
      dirty_0_210 <= _GEN_10033;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_211 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_211 <= _GEN_10034;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_211 <= _GEN_10552;
    end else begin
      dirty_0_211 <= _GEN_10034;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_212 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_212 <= _GEN_10035;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_212 <= _GEN_10553;
    end else begin
      dirty_0_212 <= _GEN_10035;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_213 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_213 <= _GEN_10036;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_213 <= _GEN_10554;
    end else begin
      dirty_0_213 <= _GEN_10036;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_214 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_214 <= _GEN_10037;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_214 <= _GEN_10555;
    end else begin
      dirty_0_214 <= _GEN_10037;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_215 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_215 <= _GEN_10038;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_215 <= _GEN_10556;
    end else begin
      dirty_0_215 <= _GEN_10038;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_216 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_216 <= _GEN_10039;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_216 <= _GEN_10557;
    end else begin
      dirty_0_216 <= _GEN_10039;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_217 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_217 <= _GEN_10040;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_217 <= _GEN_10558;
    end else begin
      dirty_0_217 <= _GEN_10040;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_218 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_218 <= _GEN_10041;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_218 <= _GEN_10559;
    end else begin
      dirty_0_218 <= _GEN_10041;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_219 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_219 <= _GEN_10042;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_219 <= _GEN_10560;
    end else begin
      dirty_0_219 <= _GEN_10042;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_220 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_220 <= _GEN_10043;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_220 <= _GEN_10561;
    end else begin
      dirty_0_220 <= _GEN_10043;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_221 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_221 <= _GEN_10044;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_221 <= _GEN_10562;
    end else begin
      dirty_0_221 <= _GEN_10044;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_222 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_222 <= _GEN_10045;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_222 <= _GEN_10563;
    end else begin
      dirty_0_222 <= _GEN_10045;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_223 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_223 <= _GEN_10046;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_223 <= _GEN_10564;
    end else begin
      dirty_0_223 <= _GEN_10046;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_224 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_224 <= _GEN_10047;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_224 <= _GEN_10565;
    end else begin
      dirty_0_224 <= _GEN_10047;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_225 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_225 <= _GEN_10048;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_225 <= _GEN_10566;
    end else begin
      dirty_0_225 <= _GEN_10048;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_226 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_226 <= _GEN_10049;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_226 <= _GEN_10567;
    end else begin
      dirty_0_226 <= _GEN_10049;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_227 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_227 <= _GEN_10050;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_227 <= _GEN_10568;
    end else begin
      dirty_0_227 <= _GEN_10050;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_228 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_228 <= _GEN_10051;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_228 <= _GEN_10569;
    end else begin
      dirty_0_228 <= _GEN_10051;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_229 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_229 <= _GEN_10052;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_229 <= _GEN_10570;
    end else begin
      dirty_0_229 <= _GEN_10052;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_230 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_230 <= _GEN_10053;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_230 <= _GEN_10571;
    end else begin
      dirty_0_230 <= _GEN_10053;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_231 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_231 <= _GEN_10054;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_231 <= _GEN_10572;
    end else begin
      dirty_0_231 <= _GEN_10054;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_232 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_232 <= _GEN_10055;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_232 <= _GEN_10573;
    end else begin
      dirty_0_232 <= _GEN_10055;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_233 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_233 <= _GEN_10056;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_233 <= _GEN_10574;
    end else begin
      dirty_0_233 <= _GEN_10056;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_234 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_234 <= _GEN_10057;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_234 <= _GEN_10575;
    end else begin
      dirty_0_234 <= _GEN_10057;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_235 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_235 <= _GEN_10058;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_235 <= _GEN_10576;
    end else begin
      dirty_0_235 <= _GEN_10058;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_236 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_236 <= _GEN_10059;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_236 <= _GEN_10577;
    end else begin
      dirty_0_236 <= _GEN_10059;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_237 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_237 <= _GEN_10060;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_237 <= _GEN_10578;
    end else begin
      dirty_0_237 <= _GEN_10060;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_238 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_238 <= _GEN_10061;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_238 <= _GEN_10579;
    end else begin
      dirty_0_238 <= _GEN_10061;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_239 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_239 <= _GEN_10062;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_239 <= _GEN_10580;
    end else begin
      dirty_0_239 <= _GEN_10062;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_240 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_240 <= _GEN_10063;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_240 <= _GEN_10581;
    end else begin
      dirty_0_240 <= _GEN_10063;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_241 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_241 <= _GEN_10064;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_241 <= _GEN_10582;
    end else begin
      dirty_0_241 <= _GEN_10064;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_242 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_242 <= _GEN_10065;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_242 <= _GEN_10583;
    end else begin
      dirty_0_242 <= _GEN_10065;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_243 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_243 <= _GEN_10066;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_243 <= _GEN_10584;
    end else begin
      dirty_0_243 <= _GEN_10066;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_244 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_244 <= _GEN_10067;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_244 <= _GEN_10585;
    end else begin
      dirty_0_244 <= _GEN_10067;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_245 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_245 <= _GEN_10068;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_245 <= _GEN_10586;
    end else begin
      dirty_0_245 <= _GEN_10068;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_246 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_246 <= _GEN_10069;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_246 <= _GEN_10587;
    end else begin
      dirty_0_246 <= _GEN_10069;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_247 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_247 <= _GEN_10070;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_247 <= _GEN_10588;
    end else begin
      dirty_0_247 <= _GEN_10070;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_248 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_248 <= _GEN_10071;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_248 <= _GEN_10589;
    end else begin
      dirty_0_248 <= _GEN_10071;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_249 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_249 <= _GEN_10072;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_249 <= _GEN_10590;
    end else begin
      dirty_0_249 <= _GEN_10072;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_250 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_250 <= _GEN_10073;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_250 <= _GEN_10591;
    end else begin
      dirty_0_250 <= _GEN_10073;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_251 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_251 <= _GEN_10074;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_251 <= _GEN_10592;
    end else begin
      dirty_0_251 <= _GEN_10074;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_252 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_252 <= _GEN_10075;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_252 <= _GEN_10593;
    end else begin
      dirty_0_252 <= _GEN_10075;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_253 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_253 <= _GEN_10076;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_253 <= _GEN_10594;
    end else begin
      dirty_0_253 <= _GEN_10076;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_254 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_254 <= _GEN_10077;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_254 <= _GEN_10595;
    end else begin
      dirty_0_254 <= _GEN_10077;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_0_255 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_255 <= _GEN_10078;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_0_255 <= _GEN_10596;
    end else begin
      dirty_0_255 <= _GEN_10078;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_0 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_0 <= _GEN_10079;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_0 <= _GEN_10597;
    end else begin
      dirty_1_0 <= _GEN_10079;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_1 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_1 <= _GEN_10080;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_1 <= _GEN_10598;
    end else begin
      dirty_1_1 <= _GEN_10080;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_2 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_2 <= _GEN_10081;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_2 <= _GEN_10599;
    end else begin
      dirty_1_2 <= _GEN_10081;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_3 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_3 <= _GEN_10082;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_3 <= _GEN_10600;
    end else begin
      dirty_1_3 <= _GEN_10082;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_4 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_4 <= _GEN_10083;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_4 <= _GEN_10601;
    end else begin
      dirty_1_4 <= _GEN_10083;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_5 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_5 <= _GEN_10084;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_5 <= _GEN_10602;
    end else begin
      dirty_1_5 <= _GEN_10084;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_6 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_6 <= _GEN_10085;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_6 <= _GEN_10603;
    end else begin
      dirty_1_6 <= _GEN_10085;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_7 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_7 <= _GEN_10086;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_7 <= _GEN_10604;
    end else begin
      dirty_1_7 <= _GEN_10086;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_8 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_8 <= _GEN_10087;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_8 <= _GEN_10605;
    end else begin
      dirty_1_8 <= _GEN_10087;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_9 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_9 <= _GEN_10088;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_9 <= _GEN_10606;
    end else begin
      dirty_1_9 <= _GEN_10088;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_10 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_10 <= _GEN_10089;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_10 <= _GEN_10607;
    end else begin
      dirty_1_10 <= _GEN_10089;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_11 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_11 <= _GEN_10090;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_11 <= _GEN_10608;
    end else begin
      dirty_1_11 <= _GEN_10090;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_12 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_12 <= _GEN_10091;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_12 <= _GEN_10609;
    end else begin
      dirty_1_12 <= _GEN_10091;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_13 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_13 <= _GEN_10092;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_13 <= _GEN_10610;
    end else begin
      dirty_1_13 <= _GEN_10092;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_14 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_14 <= _GEN_10093;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_14 <= _GEN_10611;
    end else begin
      dirty_1_14 <= _GEN_10093;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_15 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_15 <= _GEN_10094;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_15 <= _GEN_10612;
    end else begin
      dirty_1_15 <= _GEN_10094;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_16 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_16 <= _GEN_10095;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_16 <= _GEN_10613;
    end else begin
      dirty_1_16 <= _GEN_10095;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_17 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_17 <= _GEN_10096;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_17 <= _GEN_10614;
    end else begin
      dirty_1_17 <= _GEN_10096;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_18 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_18 <= _GEN_10097;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_18 <= _GEN_10615;
    end else begin
      dirty_1_18 <= _GEN_10097;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_19 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_19 <= _GEN_10098;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_19 <= _GEN_10616;
    end else begin
      dirty_1_19 <= _GEN_10098;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_20 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_20 <= _GEN_10099;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_20 <= _GEN_10617;
    end else begin
      dirty_1_20 <= _GEN_10099;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_21 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_21 <= _GEN_10100;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_21 <= _GEN_10618;
    end else begin
      dirty_1_21 <= _GEN_10100;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_22 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_22 <= _GEN_10101;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_22 <= _GEN_10619;
    end else begin
      dirty_1_22 <= _GEN_10101;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_23 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_23 <= _GEN_10102;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_23 <= _GEN_10620;
    end else begin
      dirty_1_23 <= _GEN_10102;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_24 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_24 <= _GEN_10103;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_24 <= _GEN_10621;
    end else begin
      dirty_1_24 <= _GEN_10103;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_25 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_25 <= _GEN_10104;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_25 <= _GEN_10622;
    end else begin
      dirty_1_25 <= _GEN_10104;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_26 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_26 <= _GEN_10105;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_26 <= _GEN_10623;
    end else begin
      dirty_1_26 <= _GEN_10105;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_27 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_27 <= _GEN_10106;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_27 <= _GEN_10624;
    end else begin
      dirty_1_27 <= _GEN_10106;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_28 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_28 <= _GEN_10107;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_28 <= _GEN_10625;
    end else begin
      dirty_1_28 <= _GEN_10107;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_29 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_29 <= _GEN_10108;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_29 <= _GEN_10626;
    end else begin
      dirty_1_29 <= _GEN_10108;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_30 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_30 <= _GEN_10109;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_30 <= _GEN_10627;
    end else begin
      dirty_1_30 <= _GEN_10109;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_31 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_31 <= _GEN_10110;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_31 <= _GEN_10628;
    end else begin
      dirty_1_31 <= _GEN_10110;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_32 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_32 <= _GEN_10111;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_32 <= _GEN_10629;
    end else begin
      dirty_1_32 <= _GEN_10111;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_33 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_33 <= _GEN_10112;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_33 <= _GEN_10630;
    end else begin
      dirty_1_33 <= _GEN_10112;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_34 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_34 <= _GEN_10113;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_34 <= _GEN_10631;
    end else begin
      dirty_1_34 <= _GEN_10113;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_35 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_35 <= _GEN_10114;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_35 <= _GEN_10632;
    end else begin
      dirty_1_35 <= _GEN_10114;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_36 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_36 <= _GEN_10115;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_36 <= _GEN_10633;
    end else begin
      dirty_1_36 <= _GEN_10115;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_37 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_37 <= _GEN_10116;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_37 <= _GEN_10634;
    end else begin
      dirty_1_37 <= _GEN_10116;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_38 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_38 <= _GEN_10117;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_38 <= _GEN_10635;
    end else begin
      dirty_1_38 <= _GEN_10117;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_39 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_39 <= _GEN_10118;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_39 <= _GEN_10636;
    end else begin
      dirty_1_39 <= _GEN_10118;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_40 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_40 <= _GEN_10119;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_40 <= _GEN_10637;
    end else begin
      dirty_1_40 <= _GEN_10119;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_41 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_41 <= _GEN_10120;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_41 <= _GEN_10638;
    end else begin
      dirty_1_41 <= _GEN_10120;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_42 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_42 <= _GEN_10121;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_42 <= _GEN_10639;
    end else begin
      dirty_1_42 <= _GEN_10121;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_43 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_43 <= _GEN_10122;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_43 <= _GEN_10640;
    end else begin
      dirty_1_43 <= _GEN_10122;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_44 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_44 <= _GEN_10123;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_44 <= _GEN_10641;
    end else begin
      dirty_1_44 <= _GEN_10123;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_45 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_45 <= _GEN_10124;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_45 <= _GEN_10642;
    end else begin
      dirty_1_45 <= _GEN_10124;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_46 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_46 <= _GEN_10125;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_46 <= _GEN_10643;
    end else begin
      dirty_1_46 <= _GEN_10125;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_47 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_47 <= _GEN_10126;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_47 <= _GEN_10644;
    end else begin
      dirty_1_47 <= _GEN_10126;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_48 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_48 <= _GEN_10127;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_48 <= _GEN_10645;
    end else begin
      dirty_1_48 <= _GEN_10127;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_49 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_49 <= _GEN_10128;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_49 <= _GEN_10646;
    end else begin
      dirty_1_49 <= _GEN_10128;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_50 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_50 <= _GEN_10129;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_50 <= _GEN_10647;
    end else begin
      dirty_1_50 <= _GEN_10129;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_51 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_51 <= _GEN_10130;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_51 <= _GEN_10648;
    end else begin
      dirty_1_51 <= _GEN_10130;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_52 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_52 <= _GEN_10131;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_52 <= _GEN_10649;
    end else begin
      dirty_1_52 <= _GEN_10131;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_53 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_53 <= _GEN_10132;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_53 <= _GEN_10650;
    end else begin
      dirty_1_53 <= _GEN_10132;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_54 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_54 <= _GEN_10133;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_54 <= _GEN_10651;
    end else begin
      dirty_1_54 <= _GEN_10133;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_55 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_55 <= _GEN_10134;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_55 <= _GEN_10652;
    end else begin
      dirty_1_55 <= _GEN_10134;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_56 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_56 <= _GEN_10135;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_56 <= _GEN_10653;
    end else begin
      dirty_1_56 <= _GEN_10135;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_57 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_57 <= _GEN_10136;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_57 <= _GEN_10654;
    end else begin
      dirty_1_57 <= _GEN_10136;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_58 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_58 <= _GEN_10137;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_58 <= _GEN_10655;
    end else begin
      dirty_1_58 <= _GEN_10137;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_59 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_59 <= _GEN_10138;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_59 <= _GEN_10656;
    end else begin
      dirty_1_59 <= _GEN_10138;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_60 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_60 <= _GEN_10139;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_60 <= _GEN_10657;
    end else begin
      dirty_1_60 <= _GEN_10139;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_61 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_61 <= _GEN_10140;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_61 <= _GEN_10658;
    end else begin
      dirty_1_61 <= _GEN_10140;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_62 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_62 <= _GEN_10141;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_62 <= _GEN_10659;
    end else begin
      dirty_1_62 <= _GEN_10141;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_63 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_63 <= _GEN_10142;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_63 <= _GEN_10660;
    end else begin
      dirty_1_63 <= _GEN_10142;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_64 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_64 <= _GEN_10143;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_64 <= _GEN_10661;
    end else begin
      dirty_1_64 <= _GEN_10143;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_65 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_65 <= _GEN_10144;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_65 <= _GEN_10662;
    end else begin
      dirty_1_65 <= _GEN_10144;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_66 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_66 <= _GEN_10145;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_66 <= _GEN_10663;
    end else begin
      dirty_1_66 <= _GEN_10145;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_67 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_67 <= _GEN_10146;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_67 <= _GEN_10664;
    end else begin
      dirty_1_67 <= _GEN_10146;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_68 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_68 <= _GEN_10147;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_68 <= _GEN_10665;
    end else begin
      dirty_1_68 <= _GEN_10147;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_69 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_69 <= _GEN_10148;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_69 <= _GEN_10666;
    end else begin
      dirty_1_69 <= _GEN_10148;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_70 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_70 <= _GEN_10149;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_70 <= _GEN_10667;
    end else begin
      dirty_1_70 <= _GEN_10149;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_71 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_71 <= _GEN_10150;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_71 <= _GEN_10668;
    end else begin
      dirty_1_71 <= _GEN_10150;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_72 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_72 <= _GEN_10151;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_72 <= _GEN_10669;
    end else begin
      dirty_1_72 <= _GEN_10151;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_73 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_73 <= _GEN_10152;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_73 <= _GEN_10670;
    end else begin
      dirty_1_73 <= _GEN_10152;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_74 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_74 <= _GEN_10153;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_74 <= _GEN_10671;
    end else begin
      dirty_1_74 <= _GEN_10153;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_75 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_75 <= _GEN_10154;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_75 <= _GEN_10672;
    end else begin
      dirty_1_75 <= _GEN_10154;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_76 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_76 <= _GEN_10155;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_76 <= _GEN_10673;
    end else begin
      dirty_1_76 <= _GEN_10155;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_77 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_77 <= _GEN_10156;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_77 <= _GEN_10674;
    end else begin
      dirty_1_77 <= _GEN_10156;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_78 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_78 <= _GEN_10157;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_78 <= _GEN_10675;
    end else begin
      dirty_1_78 <= _GEN_10157;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_79 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_79 <= _GEN_10158;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_79 <= _GEN_10676;
    end else begin
      dirty_1_79 <= _GEN_10158;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_80 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_80 <= _GEN_10159;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_80 <= _GEN_10677;
    end else begin
      dirty_1_80 <= _GEN_10159;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_81 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_81 <= _GEN_10160;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_81 <= _GEN_10678;
    end else begin
      dirty_1_81 <= _GEN_10160;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_82 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_82 <= _GEN_10161;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_82 <= _GEN_10679;
    end else begin
      dirty_1_82 <= _GEN_10161;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_83 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_83 <= _GEN_10162;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_83 <= _GEN_10680;
    end else begin
      dirty_1_83 <= _GEN_10162;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_84 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_84 <= _GEN_10163;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_84 <= _GEN_10681;
    end else begin
      dirty_1_84 <= _GEN_10163;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_85 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_85 <= _GEN_10164;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_85 <= _GEN_10682;
    end else begin
      dirty_1_85 <= _GEN_10164;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_86 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_86 <= _GEN_10165;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_86 <= _GEN_10683;
    end else begin
      dirty_1_86 <= _GEN_10165;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_87 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_87 <= _GEN_10166;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_87 <= _GEN_10684;
    end else begin
      dirty_1_87 <= _GEN_10166;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_88 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_88 <= _GEN_10167;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_88 <= _GEN_10685;
    end else begin
      dirty_1_88 <= _GEN_10167;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_89 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_89 <= _GEN_10168;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_89 <= _GEN_10686;
    end else begin
      dirty_1_89 <= _GEN_10168;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_90 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_90 <= _GEN_10169;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_90 <= _GEN_10687;
    end else begin
      dirty_1_90 <= _GEN_10169;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_91 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_91 <= _GEN_10170;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_91 <= _GEN_10688;
    end else begin
      dirty_1_91 <= _GEN_10170;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_92 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_92 <= _GEN_10171;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_92 <= _GEN_10689;
    end else begin
      dirty_1_92 <= _GEN_10171;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_93 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_93 <= _GEN_10172;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_93 <= _GEN_10690;
    end else begin
      dirty_1_93 <= _GEN_10172;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_94 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_94 <= _GEN_10173;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_94 <= _GEN_10691;
    end else begin
      dirty_1_94 <= _GEN_10173;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_95 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_95 <= _GEN_10174;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_95 <= _GEN_10692;
    end else begin
      dirty_1_95 <= _GEN_10174;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_96 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_96 <= _GEN_10175;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_96 <= _GEN_10693;
    end else begin
      dirty_1_96 <= _GEN_10175;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_97 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_97 <= _GEN_10176;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_97 <= _GEN_10694;
    end else begin
      dirty_1_97 <= _GEN_10176;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_98 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_98 <= _GEN_10177;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_98 <= _GEN_10695;
    end else begin
      dirty_1_98 <= _GEN_10177;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_99 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_99 <= _GEN_10178;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_99 <= _GEN_10696;
    end else begin
      dirty_1_99 <= _GEN_10178;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_100 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_100 <= _GEN_10179;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_100 <= _GEN_10697;
    end else begin
      dirty_1_100 <= _GEN_10179;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_101 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_101 <= _GEN_10180;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_101 <= _GEN_10698;
    end else begin
      dirty_1_101 <= _GEN_10180;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_102 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_102 <= _GEN_10181;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_102 <= _GEN_10699;
    end else begin
      dirty_1_102 <= _GEN_10181;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_103 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_103 <= _GEN_10182;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_103 <= _GEN_10700;
    end else begin
      dirty_1_103 <= _GEN_10182;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_104 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_104 <= _GEN_10183;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_104 <= _GEN_10701;
    end else begin
      dirty_1_104 <= _GEN_10183;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_105 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_105 <= _GEN_10184;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_105 <= _GEN_10702;
    end else begin
      dirty_1_105 <= _GEN_10184;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_106 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_106 <= _GEN_10185;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_106 <= _GEN_10703;
    end else begin
      dirty_1_106 <= _GEN_10185;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_107 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_107 <= _GEN_10186;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_107 <= _GEN_10704;
    end else begin
      dirty_1_107 <= _GEN_10186;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_108 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_108 <= _GEN_10187;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_108 <= _GEN_10705;
    end else begin
      dirty_1_108 <= _GEN_10187;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_109 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_109 <= _GEN_10188;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_109 <= _GEN_10706;
    end else begin
      dirty_1_109 <= _GEN_10188;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_110 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_110 <= _GEN_10189;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_110 <= _GEN_10707;
    end else begin
      dirty_1_110 <= _GEN_10189;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_111 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_111 <= _GEN_10190;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_111 <= _GEN_10708;
    end else begin
      dirty_1_111 <= _GEN_10190;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_112 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_112 <= _GEN_10191;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_112 <= _GEN_10709;
    end else begin
      dirty_1_112 <= _GEN_10191;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_113 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_113 <= _GEN_10192;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_113 <= _GEN_10710;
    end else begin
      dirty_1_113 <= _GEN_10192;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_114 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_114 <= _GEN_10193;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_114 <= _GEN_10711;
    end else begin
      dirty_1_114 <= _GEN_10193;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_115 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_115 <= _GEN_10194;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_115 <= _GEN_10712;
    end else begin
      dirty_1_115 <= _GEN_10194;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_116 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_116 <= _GEN_10195;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_116 <= _GEN_10713;
    end else begin
      dirty_1_116 <= _GEN_10195;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_117 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_117 <= _GEN_10196;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_117 <= _GEN_10714;
    end else begin
      dirty_1_117 <= _GEN_10196;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_118 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_118 <= _GEN_10197;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_118 <= _GEN_10715;
    end else begin
      dirty_1_118 <= _GEN_10197;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_119 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_119 <= _GEN_10198;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_119 <= _GEN_10716;
    end else begin
      dirty_1_119 <= _GEN_10198;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_120 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_120 <= _GEN_10199;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_120 <= _GEN_10717;
    end else begin
      dirty_1_120 <= _GEN_10199;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_121 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_121 <= _GEN_10200;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_121 <= _GEN_10718;
    end else begin
      dirty_1_121 <= _GEN_10200;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_122 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_122 <= _GEN_10201;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_122 <= _GEN_10719;
    end else begin
      dirty_1_122 <= _GEN_10201;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_123 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_123 <= _GEN_10202;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_123 <= _GEN_10720;
    end else begin
      dirty_1_123 <= _GEN_10202;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_124 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_124 <= _GEN_10203;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_124 <= _GEN_10721;
    end else begin
      dirty_1_124 <= _GEN_10203;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_125 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_125 <= _GEN_10204;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_125 <= _GEN_10722;
    end else begin
      dirty_1_125 <= _GEN_10204;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_126 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_126 <= _GEN_10205;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_126 <= _GEN_10723;
    end else begin
      dirty_1_126 <= _GEN_10205;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_127 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_127 <= _GEN_10206;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_127 <= _GEN_10724;
    end else begin
      dirty_1_127 <= _GEN_10206;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_128 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_128 <= _GEN_10207;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_128 <= _GEN_10725;
    end else begin
      dirty_1_128 <= _GEN_10207;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_129 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_129 <= _GEN_10208;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_129 <= _GEN_10726;
    end else begin
      dirty_1_129 <= _GEN_10208;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_130 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_130 <= _GEN_10209;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_130 <= _GEN_10727;
    end else begin
      dirty_1_130 <= _GEN_10209;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_131 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_131 <= _GEN_10210;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_131 <= _GEN_10728;
    end else begin
      dirty_1_131 <= _GEN_10210;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_132 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_132 <= _GEN_10211;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_132 <= _GEN_10729;
    end else begin
      dirty_1_132 <= _GEN_10211;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_133 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_133 <= _GEN_10212;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_133 <= _GEN_10730;
    end else begin
      dirty_1_133 <= _GEN_10212;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_134 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_134 <= _GEN_10213;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_134 <= _GEN_10731;
    end else begin
      dirty_1_134 <= _GEN_10213;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_135 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_135 <= _GEN_10214;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_135 <= _GEN_10732;
    end else begin
      dirty_1_135 <= _GEN_10214;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_136 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_136 <= _GEN_10215;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_136 <= _GEN_10733;
    end else begin
      dirty_1_136 <= _GEN_10215;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_137 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_137 <= _GEN_10216;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_137 <= _GEN_10734;
    end else begin
      dirty_1_137 <= _GEN_10216;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_138 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_138 <= _GEN_10217;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_138 <= _GEN_10735;
    end else begin
      dirty_1_138 <= _GEN_10217;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_139 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_139 <= _GEN_10218;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_139 <= _GEN_10736;
    end else begin
      dirty_1_139 <= _GEN_10218;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_140 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_140 <= _GEN_10219;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_140 <= _GEN_10737;
    end else begin
      dirty_1_140 <= _GEN_10219;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_141 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_141 <= _GEN_10220;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_141 <= _GEN_10738;
    end else begin
      dirty_1_141 <= _GEN_10220;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_142 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_142 <= _GEN_10221;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_142 <= _GEN_10739;
    end else begin
      dirty_1_142 <= _GEN_10221;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_143 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_143 <= _GEN_10222;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_143 <= _GEN_10740;
    end else begin
      dirty_1_143 <= _GEN_10222;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_144 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_144 <= _GEN_10223;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_144 <= _GEN_10741;
    end else begin
      dirty_1_144 <= _GEN_10223;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_145 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_145 <= _GEN_10224;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_145 <= _GEN_10742;
    end else begin
      dirty_1_145 <= _GEN_10224;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_146 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_146 <= _GEN_10225;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_146 <= _GEN_10743;
    end else begin
      dirty_1_146 <= _GEN_10225;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_147 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_147 <= _GEN_10226;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_147 <= _GEN_10744;
    end else begin
      dirty_1_147 <= _GEN_10226;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_148 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_148 <= _GEN_10227;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_148 <= _GEN_10745;
    end else begin
      dirty_1_148 <= _GEN_10227;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_149 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_149 <= _GEN_10228;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_149 <= _GEN_10746;
    end else begin
      dirty_1_149 <= _GEN_10228;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_150 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_150 <= _GEN_10229;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_150 <= _GEN_10747;
    end else begin
      dirty_1_150 <= _GEN_10229;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_151 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_151 <= _GEN_10230;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_151 <= _GEN_10748;
    end else begin
      dirty_1_151 <= _GEN_10230;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_152 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_152 <= _GEN_10231;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_152 <= _GEN_10749;
    end else begin
      dirty_1_152 <= _GEN_10231;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_153 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_153 <= _GEN_10232;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_153 <= _GEN_10750;
    end else begin
      dirty_1_153 <= _GEN_10232;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_154 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_154 <= _GEN_10233;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_154 <= _GEN_10751;
    end else begin
      dirty_1_154 <= _GEN_10233;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_155 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_155 <= _GEN_10234;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_155 <= _GEN_10752;
    end else begin
      dirty_1_155 <= _GEN_10234;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_156 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_156 <= _GEN_10235;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_156 <= _GEN_10753;
    end else begin
      dirty_1_156 <= _GEN_10235;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_157 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_157 <= _GEN_10236;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_157 <= _GEN_10754;
    end else begin
      dirty_1_157 <= _GEN_10236;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_158 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_158 <= _GEN_10237;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_158 <= _GEN_10755;
    end else begin
      dirty_1_158 <= _GEN_10237;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_159 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_159 <= _GEN_10238;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_159 <= _GEN_10756;
    end else begin
      dirty_1_159 <= _GEN_10238;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_160 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_160 <= _GEN_10239;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_160 <= _GEN_10757;
    end else begin
      dirty_1_160 <= _GEN_10239;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_161 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_161 <= _GEN_10240;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_161 <= _GEN_10758;
    end else begin
      dirty_1_161 <= _GEN_10240;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_162 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_162 <= _GEN_10241;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_162 <= _GEN_10759;
    end else begin
      dirty_1_162 <= _GEN_10241;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_163 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_163 <= _GEN_10242;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_163 <= _GEN_10760;
    end else begin
      dirty_1_163 <= _GEN_10242;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_164 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_164 <= _GEN_10243;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_164 <= _GEN_10761;
    end else begin
      dirty_1_164 <= _GEN_10243;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_165 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_165 <= _GEN_10244;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_165 <= _GEN_10762;
    end else begin
      dirty_1_165 <= _GEN_10244;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_166 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_166 <= _GEN_10245;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_166 <= _GEN_10763;
    end else begin
      dirty_1_166 <= _GEN_10245;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_167 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_167 <= _GEN_10246;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_167 <= _GEN_10764;
    end else begin
      dirty_1_167 <= _GEN_10246;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_168 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_168 <= _GEN_10247;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_168 <= _GEN_10765;
    end else begin
      dirty_1_168 <= _GEN_10247;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_169 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_169 <= _GEN_10248;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_169 <= _GEN_10766;
    end else begin
      dirty_1_169 <= _GEN_10248;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_170 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_170 <= _GEN_10249;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_170 <= _GEN_10767;
    end else begin
      dirty_1_170 <= _GEN_10249;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_171 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_171 <= _GEN_10250;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_171 <= _GEN_10768;
    end else begin
      dirty_1_171 <= _GEN_10250;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_172 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_172 <= _GEN_10251;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_172 <= _GEN_10769;
    end else begin
      dirty_1_172 <= _GEN_10251;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_173 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_173 <= _GEN_10252;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_173 <= _GEN_10770;
    end else begin
      dirty_1_173 <= _GEN_10252;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_174 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_174 <= _GEN_10253;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_174 <= _GEN_10771;
    end else begin
      dirty_1_174 <= _GEN_10253;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_175 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_175 <= _GEN_10254;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_175 <= _GEN_10772;
    end else begin
      dirty_1_175 <= _GEN_10254;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_176 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_176 <= _GEN_10255;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_176 <= _GEN_10773;
    end else begin
      dirty_1_176 <= _GEN_10255;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_177 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_177 <= _GEN_10256;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_177 <= _GEN_10774;
    end else begin
      dirty_1_177 <= _GEN_10256;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_178 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_178 <= _GEN_10257;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_178 <= _GEN_10775;
    end else begin
      dirty_1_178 <= _GEN_10257;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_179 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_179 <= _GEN_10258;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_179 <= _GEN_10776;
    end else begin
      dirty_1_179 <= _GEN_10258;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_180 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_180 <= _GEN_10259;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_180 <= _GEN_10777;
    end else begin
      dirty_1_180 <= _GEN_10259;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_181 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_181 <= _GEN_10260;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_181 <= _GEN_10778;
    end else begin
      dirty_1_181 <= _GEN_10260;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_182 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_182 <= _GEN_10261;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_182 <= _GEN_10779;
    end else begin
      dirty_1_182 <= _GEN_10261;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_183 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_183 <= _GEN_10262;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_183 <= _GEN_10780;
    end else begin
      dirty_1_183 <= _GEN_10262;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_184 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_184 <= _GEN_10263;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_184 <= _GEN_10781;
    end else begin
      dirty_1_184 <= _GEN_10263;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_185 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_185 <= _GEN_10264;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_185 <= _GEN_10782;
    end else begin
      dirty_1_185 <= _GEN_10264;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_186 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_186 <= _GEN_10265;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_186 <= _GEN_10783;
    end else begin
      dirty_1_186 <= _GEN_10265;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_187 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_187 <= _GEN_10266;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_187 <= _GEN_10784;
    end else begin
      dirty_1_187 <= _GEN_10266;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_188 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_188 <= _GEN_10267;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_188 <= _GEN_10785;
    end else begin
      dirty_1_188 <= _GEN_10267;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_189 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_189 <= _GEN_10268;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_189 <= _GEN_10786;
    end else begin
      dirty_1_189 <= _GEN_10268;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_190 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_190 <= _GEN_10269;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_190 <= _GEN_10787;
    end else begin
      dirty_1_190 <= _GEN_10269;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_191 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_191 <= _GEN_10270;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_191 <= _GEN_10788;
    end else begin
      dirty_1_191 <= _GEN_10270;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_192 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_192 <= _GEN_10271;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_192 <= _GEN_10789;
    end else begin
      dirty_1_192 <= _GEN_10271;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_193 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_193 <= _GEN_10272;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_193 <= _GEN_10790;
    end else begin
      dirty_1_193 <= _GEN_10272;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_194 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_194 <= _GEN_10273;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_194 <= _GEN_10791;
    end else begin
      dirty_1_194 <= _GEN_10273;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_195 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_195 <= _GEN_10274;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_195 <= _GEN_10792;
    end else begin
      dirty_1_195 <= _GEN_10274;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_196 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_196 <= _GEN_10275;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_196 <= _GEN_10793;
    end else begin
      dirty_1_196 <= _GEN_10275;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_197 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_197 <= _GEN_10276;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_197 <= _GEN_10794;
    end else begin
      dirty_1_197 <= _GEN_10276;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_198 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_198 <= _GEN_10277;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_198 <= _GEN_10795;
    end else begin
      dirty_1_198 <= _GEN_10277;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_199 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_199 <= _GEN_10278;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_199 <= _GEN_10796;
    end else begin
      dirty_1_199 <= _GEN_10278;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_200 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_200 <= _GEN_10279;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_200 <= _GEN_10797;
    end else begin
      dirty_1_200 <= _GEN_10279;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_201 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_201 <= _GEN_10280;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_201 <= _GEN_10798;
    end else begin
      dirty_1_201 <= _GEN_10280;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_202 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_202 <= _GEN_10281;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_202 <= _GEN_10799;
    end else begin
      dirty_1_202 <= _GEN_10281;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_203 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_203 <= _GEN_10282;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_203 <= _GEN_10800;
    end else begin
      dirty_1_203 <= _GEN_10282;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_204 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_204 <= _GEN_10283;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_204 <= _GEN_10801;
    end else begin
      dirty_1_204 <= _GEN_10283;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_205 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_205 <= _GEN_10284;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_205 <= _GEN_10802;
    end else begin
      dirty_1_205 <= _GEN_10284;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_206 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_206 <= _GEN_10285;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_206 <= _GEN_10803;
    end else begin
      dirty_1_206 <= _GEN_10285;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_207 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_207 <= _GEN_10286;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_207 <= _GEN_10804;
    end else begin
      dirty_1_207 <= _GEN_10286;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_208 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_208 <= _GEN_10287;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_208 <= _GEN_10805;
    end else begin
      dirty_1_208 <= _GEN_10287;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_209 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_209 <= _GEN_10288;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_209 <= _GEN_10806;
    end else begin
      dirty_1_209 <= _GEN_10288;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_210 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_210 <= _GEN_10289;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_210 <= _GEN_10807;
    end else begin
      dirty_1_210 <= _GEN_10289;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_211 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_211 <= _GEN_10290;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_211 <= _GEN_10808;
    end else begin
      dirty_1_211 <= _GEN_10290;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_212 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_212 <= _GEN_10291;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_212 <= _GEN_10809;
    end else begin
      dirty_1_212 <= _GEN_10291;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_213 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_213 <= _GEN_10292;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_213 <= _GEN_10810;
    end else begin
      dirty_1_213 <= _GEN_10292;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_214 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_214 <= _GEN_10293;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_214 <= _GEN_10811;
    end else begin
      dirty_1_214 <= _GEN_10293;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_215 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_215 <= _GEN_10294;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_215 <= _GEN_10812;
    end else begin
      dirty_1_215 <= _GEN_10294;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_216 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_216 <= _GEN_10295;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_216 <= _GEN_10813;
    end else begin
      dirty_1_216 <= _GEN_10295;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_217 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_217 <= _GEN_10296;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_217 <= _GEN_10814;
    end else begin
      dirty_1_217 <= _GEN_10296;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_218 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_218 <= _GEN_10297;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_218 <= _GEN_10815;
    end else begin
      dirty_1_218 <= _GEN_10297;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_219 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_219 <= _GEN_10298;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_219 <= _GEN_10816;
    end else begin
      dirty_1_219 <= _GEN_10298;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_220 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_220 <= _GEN_10299;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_220 <= _GEN_10817;
    end else begin
      dirty_1_220 <= _GEN_10299;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_221 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_221 <= _GEN_10300;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_221 <= _GEN_10818;
    end else begin
      dirty_1_221 <= _GEN_10300;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_222 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_222 <= _GEN_10301;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_222 <= _GEN_10819;
    end else begin
      dirty_1_222 <= _GEN_10301;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_223 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_223 <= _GEN_10302;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_223 <= _GEN_10820;
    end else begin
      dirty_1_223 <= _GEN_10302;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_224 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_224 <= _GEN_10303;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_224 <= _GEN_10821;
    end else begin
      dirty_1_224 <= _GEN_10303;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_225 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_225 <= _GEN_10304;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_225 <= _GEN_10822;
    end else begin
      dirty_1_225 <= _GEN_10304;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_226 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_226 <= _GEN_10305;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_226 <= _GEN_10823;
    end else begin
      dirty_1_226 <= _GEN_10305;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_227 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_227 <= _GEN_10306;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_227 <= _GEN_10824;
    end else begin
      dirty_1_227 <= _GEN_10306;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_228 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_228 <= _GEN_10307;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_228 <= _GEN_10825;
    end else begin
      dirty_1_228 <= _GEN_10307;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_229 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_229 <= _GEN_10308;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_229 <= _GEN_10826;
    end else begin
      dirty_1_229 <= _GEN_10308;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_230 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_230 <= _GEN_10309;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_230 <= _GEN_10827;
    end else begin
      dirty_1_230 <= _GEN_10309;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_231 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_231 <= _GEN_10310;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_231 <= _GEN_10828;
    end else begin
      dirty_1_231 <= _GEN_10310;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_232 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_232 <= _GEN_10311;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_232 <= _GEN_10829;
    end else begin
      dirty_1_232 <= _GEN_10311;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_233 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_233 <= _GEN_10312;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_233 <= _GEN_10830;
    end else begin
      dirty_1_233 <= _GEN_10312;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_234 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_234 <= _GEN_10313;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_234 <= _GEN_10831;
    end else begin
      dirty_1_234 <= _GEN_10313;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_235 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_235 <= _GEN_10314;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_235 <= _GEN_10832;
    end else begin
      dirty_1_235 <= _GEN_10314;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_236 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_236 <= _GEN_10315;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_236 <= _GEN_10833;
    end else begin
      dirty_1_236 <= _GEN_10315;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_237 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_237 <= _GEN_10316;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_237 <= _GEN_10834;
    end else begin
      dirty_1_237 <= _GEN_10316;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_238 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_238 <= _GEN_10317;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_238 <= _GEN_10835;
    end else begin
      dirty_1_238 <= _GEN_10317;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_239 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_239 <= _GEN_10318;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_239 <= _GEN_10836;
    end else begin
      dirty_1_239 <= _GEN_10318;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_240 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_240 <= _GEN_10319;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_240 <= _GEN_10837;
    end else begin
      dirty_1_240 <= _GEN_10319;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_241 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_241 <= _GEN_10320;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_241 <= _GEN_10838;
    end else begin
      dirty_1_241 <= _GEN_10320;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_242 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_242 <= _GEN_10321;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_242 <= _GEN_10839;
    end else begin
      dirty_1_242 <= _GEN_10321;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_243 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_243 <= _GEN_10322;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_243 <= _GEN_10840;
    end else begin
      dirty_1_243 <= _GEN_10322;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_244 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_244 <= _GEN_10323;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_244 <= _GEN_10841;
    end else begin
      dirty_1_244 <= _GEN_10323;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_245 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_245 <= _GEN_10324;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_245 <= _GEN_10842;
    end else begin
      dirty_1_245 <= _GEN_10324;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_246 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_246 <= _GEN_10325;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_246 <= _GEN_10843;
    end else begin
      dirty_1_246 <= _GEN_10325;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_247 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_247 <= _GEN_10326;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_247 <= _GEN_10844;
    end else begin
      dirty_1_247 <= _GEN_10326;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_248 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_248 <= _GEN_10327;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_248 <= _GEN_10845;
    end else begin
      dirty_1_248 <= _GEN_10327;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_249 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_249 <= _GEN_10328;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_249 <= _GEN_10846;
    end else begin
      dirty_1_249 <= _GEN_10328;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_250 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_250 <= _GEN_10329;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_250 <= _GEN_10847;
    end else begin
      dirty_1_250 <= _GEN_10329;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_251 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_251 <= _GEN_10330;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_251 <= _GEN_10848;
    end else begin
      dirty_1_251 <= _GEN_10330;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_252 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_252 <= _GEN_10331;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_252 <= _GEN_10849;
    end else begin
      dirty_1_252 <= _GEN_10331;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_253 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_253 <= _GEN_10332;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_253 <= _GEN_10850;
    end else begin
      dirty_1_253 <= _GEN_10332;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_254 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_254 <= _GEN_10333;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_254 <= _GEN_10851;
    end else begin
      dirty_1_254 <= _GEN_10333;
    end
    if (reset) begin // @[dcache.scala 113:28]
      dirty_1_255 <= 1'h0; // @[dcache.scala 113:28]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_255 <= _GEN_10334;
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      dirty_1_255 <= _GEN_10852;
    end else begin
      dirty_1_255 <= _GEN_10334;
    end
    if (reset) begin // @[dcache.scala 116:34]
      req_valid <= 1'h0; // @[dcache.scala 116:34]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (!(cache_op_en)) begin // @[dcache.scala 185:30]
        if (valid) begin // @[dcache.scala 204:30]
          req_valid <= valid; // @[dcache.scala 208:33]
        end
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (!(cacheInst_r)) begin // @[dcache.scala 255:30]
        req_valid <= _GEN_114;
      end
    end else if (!(3'h2 == state)) begin // @[dcache.scala 183:18]
      req_valid <= _GEN_8626;
    end
    if (reset) begin // @[dcache.scala 118:34]
      req_op <= 1'h0; // @[dcache.scala 118:34]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        req_op <= 1'h0; // @[dcache.scala 188:33]
      end else if (valid) begin // @[dcache.scala 204:30]
        req_op <= op; // @[dcache.scala 207:33]
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (!(cacheInst_r)) begin // @[dcache.scala 255:30]
        req_op <= _GEN_117;
      end
    end
    if (reset) begin // @[dcache.scala 119:34]
      req_uncached <= 1'h0; // @[dcache.scala 119:34]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        req_uncached <= 1'h0; // @[dcache.scala 187:33]
      end else if (valid) begin // @[dcache.scala 204:30]
        req_uncached <= uncached; // @[dcache.scala 212:33]
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (!(cacheInst_r)) begin // @[dcache.scala 255:30]
        req_uncached <= _GEN_115;
      end
    end
    if (reset) begin // @[dcache.scala 120:34]
      req_offset <= 4'h0; // @[dcache.scala 120:34]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (!(cache_op_en)) begin // @[dcache.scala 185:30]
        if (valid) begin // @[dcache.scala 204:30]
          req_offset <= offset; // @[dcache.scala 211:33]
        end
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (!(cacheInst_r)) begin // @[dcache.scala 255:30]
        req_offset <= _GEN_120;
      end
    end
    if (reset) begin // @[dcache.scala 121:34]
      req_lstype <= 3'h0; // @[dcache.scala 121:34]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (!(cache_op_en)) begin // @[dcache.scala 185:30]
        if (valid) begin // @[dcache.scala 204:30]
          req_lstype <= lstype; // @[dcache.scala 213:33]
        end
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (!(cacheInst_r)) begin // @[dcache.scala 255:30]
        req_lstype <= _GEN_116;
      end
    end
    if (reset) begin // @[dcache.scala 122:34]
      req_set <= 8'h0; // @[dcache.scala 122:34]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        req_set <= cache_index; // @[dcache.scala 190:33]
      end else if (valid) begin // @[dcache.scala 204:30]
        req_set <= index; // @[dcache.scala 210:33]
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (!(cacheInst_r)) begin // @[dcache.scala 255:30]
        req_set <= _GEN_119;
      end
    end
    if (reset) begin // @[dcache.scala 123:34]
      req_tag <= 20'h0; // @[dcache.scala 123:34]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        req_tag <= cache_tag; // @[dcache.scala 189:33]
      end else if (valid) begin // @[dcache.scala 204:30]
        req_tag <= tag; // @[dcache.scala 209:33]
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (!(cacheInst_r)) begin // @[dcache.scala 255:30]
        req_tag <= _GEN_118;
      end
    end
    if (reset) begin // @[dcache.scala 124:34]
      req_wstrb_0 <= 4'h0; // @[dcache.scala 124:34]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (!(cache_op_en)) begin // @[dcache.scala 185:30]
        if (valid) begin // @[dcache.scala 204:30]
          req_wstrb_0 <= wstrb; // @[dcache.scala 214:33]
        end
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (!(cacheInst_r)) begin // @[dcache.scala 255:30]
        req_wstrb_0 <= _GEN_121;
      end
    end
    if (reset) begin // @[dcache.scala 125:34]
      req_wdata_0 <= 32'h0; // @[dcache.scala 125:34]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (!(cache_op_en)) begin // @[dcache.scala 185:30]
        if (valid) begin // @[dcache.scala 204:30]
          req_wdata_0 <= wdata; // @[dcache.scala 215:33]
        end
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (!(cacheInst_r)) begin // @[dcache.scala 255:30]
        req_wdata_0 <= _GEN_122;
      end
    end
    if (reset) begin // @[dcache.scala 127:34]
      req_wdata_1 <= 32'h0; // @[dcache.scala 127:34]
    end else if (!(3'h0 == state)) begin // @[dcache.scala 183:18]
      if (3'h1 == state) begin // @[dcache.scala 183:18]
        if (tagv_1_douta[19:0] == req_tag & tagv_1_douta[20]) begin // @[dcache.scala 226:78]
          req_wdata_1 <= _GEN_69;
        end else begin
          req_wdata_1 <= _GEN_52;
        end
      end
    end
    if (reset) begin // @[dcache.scala 128:34]
      req_wstrb_1 <= 4'h0; // @[dcache.scala 128:34]
    end else if (!(3'h0 == state)) begin // @[dcache.scala 183:18]
      if (3'h1 == state) begin // @[dcache.scala 183:18]
        if (tagv_1_douta[19:0] == req_tag & tagv_1_douta[20]) begin // @[dcache.scala 226:78]
          req_wstrb_1 <= _GEN_68;
        end else begin
          req_wstrb_1 <= _GEN_51;
        end
      end
    end
    if (reset) begin // @[dcache.scala 129:34]
      req_wline <= 1'h0; // @[dcache.scala 129:34]
    end else if (!(3'h0 == state)) begin // @[dcache.scala 183:18]
      if (3'h1 == state) begin // @[dcache.scala 183:18]
        if (tagv_1_douta[19:0] == req_tag & tagv_1_douta[20]) begin // @[dcache.scala 226:78]
          req_wline <= _GEN_67;
        end else begin
          req_wline <= _GEN_50;
        end
      end
    end
    if (reset) begin // @[dcache.scala 130:34]
      req_wset <= 8'h0; // @[dcache.scala 130:34]
    end else if (!(3'h0 == state)) begin // @[dcache.scala 183:18]
      if (3'h1 == state) begin // @[dcache.scala 183:18]
        if (tagv_1_douta[19:0] == req_tag & tagv_1_douta[20]) begin // @[dcache.scala 226:78]
          req_wset <= _GEN_66;
        end else begin
          req_wset <= _GEN_49;
        end
      end
    end
    if (reset) begin // @[dcache.scala 131:34]
      req_woffset <= 4'h0; // @[dcache.scala 131:34]
    end else if (!(3'h0 == state)) begin // @[dcache.scala 183:18]
      if (3'h1 == state) begin // @[dcache.scala 183:18]
        if (tagv_1_douta[19:0] == req_tag & tagv_1_douta[20]) begin // @[dcache.scala 226:78]
          req_woffset <= _GEN_65;
        end else begin
          req_woffset <= _GEN_48;
        end
      end
    end
    if (reset) begin // @[dcache.scala 136:34]
      tagv_r_0 <= 21'h0; // @[dcache.scala 136:34]
    end else if (!(3'h0 == state)) begin // @[dcache.scala 183:18]
      if (3'h1 == state) begin // @[dcache.scala 183:18]
        tagv_r_0 <= tagv_0_douta; // @[dcache.scala 252:29]
      end
    end
    if (reset) begin // @[dcache.scala 136:34]
      tagv_r_1 <= 21'h0; // @[dcache.scala 136:34]
    end else if (!(3'h0 == state)) begin // @[dcache.scala 183:18]
      if (3'h1 == state) begin // @[dcache.scala 183:18]
        tagv_r_1 <= tagv_1_douta; // @[dcache.scala 252:29]
      end
    end
    if (reset) begin // @[dcache.scala 171:34]
      state <= 3'h0; // @[dcache.scala 171:34]
    end else if (3'h0 == state) begin // @[dcache.scala 183:18]
      if (cache_op_en) begin // @[dcache.scala 185:30]
        state <= 3'h1; // @[dcache.scala 186:33]
      end else if (valid) begin // @[dcache.scala 204:30]
        state <= _state_T; // @[dcache.scala 205:33]
      end
    end else if (3'h1 == state) begin // @[dcache.scala 183:18]
      if (cacheInst_r) begin // @[dcache.scala 255:30]
        state <= _GEN_90;
      end else begin
        state <= _GEN_112;
      end
    end else if (3'h2 == state) begin // @[dcache.scala 183:18]
      state <= 3'h3; // @[dcache.scala 315:19]
    end else begin
      state <= _GEN_8081;
    end
    if (reset) begin // @[dcache.scala 174:34]
      refillIDX_r <= 1'h0; // @[dcache.scala 174:34]
    end else if (!(3'h0 == state)) begin // @[dcache.scala 183:18]
      if (3'h1 == state) begin // @[dcache.scala 183:18]
        if (cacheInst_r) begin // @[dcache.scala 255:30]
          refillIDX_r <= _GEN_91;
        end else begin
          refillIDX_r <= _GEN_80;
        end
      end else if (3'h2 == state) begin // @[dcache.scala 183:18]
        refillIDX_r <= refillIDX; // @[dcache.scala 331:25]
      end
    end
    LFSR_result <= {LFSR_result_hi,LFSR_result_lo}; // @[PRNG.scala 95:17]
    if (reset) begin // @[dcache.scala 178:34]
      wr_cnt <= 2'h0; // @[dcache.scala 178:34]
    end else if (!(3'h0 == state)) begin // @[dcache.scala 183:18]
      if (!(3'h1 == state)) begin // @[dcache.scala 183:18]
        if (!(3'h2 == state)) begin // @[dcache.scala 183:18]
          wr_cnt <= _GEN_8092;
        end
      end
    end
    if (reset) begin // @[dcache.scala 441:31]
      wstate <= 2'h0; // @[dcache.scala 441:31]
    end else if (2'h0 == wstate) begin // @[dcache.scala 446:19]
      if (hit & req_op) begin // @[dcache.scala 448:31]
        wstate <= 2'h1; // @[dcache.scala 449:29]
      end
    end else if (2'h1 == wstate) begin // @[dcache.scala 446:19]
      if (_T_53) begin // @[dcache.scala 460:31]
        wstate <= 2'h1; // @[dcache.scala 461:29]
      end else begin
        wstate <= 2'h2; // @[dcache.scala 464:31]
      end
    end else if (2'h2 == wstate) begin // @[dcache.scala 446:19]
      wstate <= _GEN_10878;
    end
    if (reset) begin // @[dcache.scala 444:32]
      req_wline_1 <= 1'h0; // @[dcache.scala 444:32]
    end else if (!(2'h0 == wstate)) begin // @[dcache.scala 446:19]
      if (2'h1 == wstate) begin // @[dcache.scala 446:19]
        req_wline_1 <= req_wline; // @[dcache.scala 458:61]
      end
    end
    if (reset) begin // @[dcache.scala 443:32]
      req_woffset_1 <= 4'h0; // @[dcache.scala 443:32]
    end else if (!(2'h0 == wstate)) begin // @[dcache.scala 446:19]
      if (2'h1 == wstate) begin // @[dcache.scala 446:19]
        req_woffset_1 <= req_woffset; // @[dcache.scala 459:61]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cacheInst_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  invalidate = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  loadTag = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  storeTag = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  writeBack = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  indexOnly = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dirty_0_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dirty_0_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dirty_0_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  dirty_0_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  dirty_0_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dirty_0_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  dirty_0_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  dirty_0_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dirty_0_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  dirty_0_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dirty_0_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  dirty_0_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  dirty_0_12 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  dirty_0_13 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  dirty_0_14 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  dirty_0_15 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  dirty_0_16 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  dirty_0_17 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  dirty_0_18 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  dirty_0_19 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  dirty_0_20 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  dirty_0_21 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  dirty_0_22 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  dirty_0_23 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  dirty_0_24 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  dirty_0_25 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  dirty_0_26 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  dirty_0_27 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  dirty_0_28 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  dirty_0_29 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  dirty_0_30 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  dirty_0_31 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dirty_0_32 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  dirty_0_33 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  dirty_0_34 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  dirty_0_35 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  dirty_0_36 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  dirty_0_37 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  dirty_0_38 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  dirty_0_39 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  dirty_0_40 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  dirty_0_41 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  dirty_0_42 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  dirty_0_43 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  dirty_0_44 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  dirty_0_45 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  dirty_0_46 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  dirty_0_47 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  dirty_0_48 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  dirty_0_49 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  dirty_0_50 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  dirty_0_51 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  dirty_0_52 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  dirty_0_53 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  dirty_0_54 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  dirty_0_55 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  dirty_0_56 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  dirty_0_57 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  dirty_0_58 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  dirty_0_59 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  dirty_0_60 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  dirty_0_61 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dirty_0_62 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dirty_0_63 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  dirty_0_64 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dirty_0_65 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  dirty_0_66 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  dirty_0_67 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dirty_0_68 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  dirty_0_69 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dirty_0_70 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dirty_0_71 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  dirty_0_72 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  dirty_0_73 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dirty_0_74 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  dirty_0_75 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  dirty_0_76 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  dirty_0_77 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  dirty_0_78 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  dirty_0_79 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dirty_0_80 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  dirty_0_81 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  dirty_0_82 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  dirty_0_83 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  dirty_0_84 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  dirty_0_85 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  dirty_0_86 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  dirty_0_87 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  dirty_0_88 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  dirty_0_89 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  dirty_0_90 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  dirty_0_91 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  dirty_0_92 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  dirty_0_93 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  dirty_0_94 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  dirty_0_95 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  dirty_0_96 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  dirty_0_97 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  dirty_0_98 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  dirty_0_99 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  dirty_0_100 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  dirty_0_101 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  dirty_0_102 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  dirty_0_103 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  dirty_0_104 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  dirty_0_105 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  dirty_0_106 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  dirty_0_107 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  dirty_0_108 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  dirty_0_109 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  dirty_0_110 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  dirty_0_111 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  dirty_0_112 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  dirty_0_113 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  dirty_0_114 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  dirty_0_115 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  dirty_0_116 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  dirty_0_117 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  dirty_0_118 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  dirty_0_119 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  dirty_0_120 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  dirty_0_121 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dirty_0_122 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  dirty_0_123 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  dirty_0_124 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  dirty_0_125 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  dirty_0_126 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  dirty_0_127 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  dirty_0_128 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  dirty_0_129 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  dirty_0_130 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  dirty_0_131 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  dirty_0_132 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  dirty_0_133 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  dirty_0_134 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  dirty_0_135 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  dirty_0_136 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  dirty_0_137 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  dirty_0_138 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  dirty_0_139 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  dirty_0_140 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  dirty_0_141 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  dirty_0_142 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  dirty_0_143 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  dirty_0_144 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  dirty_0_145 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  dirty_0_146 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  dirty_0_147 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  dirty_0_148 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  dirty_0_149 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  dirty_0_150 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  dirty_0_151 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  dirty_0_152 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  dirty_0_153 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  dirty_0_154 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  dirty_0_155 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  dirty_0_156 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  dirty_0_157 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  dirty_0_158 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  dirty_0_159 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  dirty_0_160 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  dirty_0_161 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  dirty_0_162 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  dirty_0_163 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  dirty_0_164 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  dirty_0_165 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  dirty_0_166 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  dirty_0_167 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  dirty_0_168 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  dirty_0_169 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  dirty_0_170 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  dirty_0_171 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  dirty_0_172 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  dirty_0_173 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  dirty_0_174 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  dirty_0_175 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  dirty_0_176 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  dirty_0_177 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  dirty_0_178 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  dirty_0_179 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  dirty_0_180 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  dirty_0_181 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  dirty_0_182 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  dirty_0_183 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  dirty_0_184 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  dirty_0_185 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  dirty_0_186 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  dirty_0_187 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  dirty_0_188 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  dirty_0_189 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  dirty_0_190 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  dirty_0_191 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  dirty_0_192 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  dirty_0_193 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  dirty_0_194 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  dirty_0_195 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  dirty_0_196 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  dirty_0_197 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  dirty_0_198 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  dirty_0_199 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  dirty_0_200 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  dirty_0_201 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  dirty_0_202 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  dirty_0_203 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  dirty_0_204 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  dirty_0_205 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dirty_0_206 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  dirty_0_207 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  dirty_0_208 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  dirty_0_209 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  dirty_0_210 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  dirty_0_211 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  dirty_0_212 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  dirty_0_213 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  dirty_0_214 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  dirty_0_215 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  dirty_0_216 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  dirty_0_217 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  dirty_0_218 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  dirty_0_219 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  dirty_0_220 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  dirty_0_221 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  dirty_0_222 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  dirty_0_223 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  dirty_0_224 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  dirty_0_225 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  dirty_0_226 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  dirty_0_227 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  dirty_0_228 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  dirty_0_229 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  dirty_0_230 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  dirty_0_231 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  dirty_0_232 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  dirty_0_233 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  dirty_0_234 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  dirty_0_235 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  dirty_0_236 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  dirty_0_237 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  dirty_0_238 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  dirty_0_239 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  dirty_0_240 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  dirty_0_241 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  dirty_0_242 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  dirty_0_243 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  dirty_0_244 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  dirty_0_245 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  dirty_0_246 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  dirty_0_247 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  dirty_0_248 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  dirty_0_249 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  dirty_0_250 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  dirty_0_251 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  dirty_0_252 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  dirty_0_253 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  dirty_0_254 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  dirty_0_255 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  dirty_1_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  dirty_1_1 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  dirty_1_2 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  dirty_1_3 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  dirty_1_4 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  dirty_1_5 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  dirty_1_6 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  dirty_1_7 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  dirty_1_8 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  dirty_1_9 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  dirty_1_10 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  dirty_1_11 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  dirty_1_12 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  dirty_1_13 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  dirty_1_14 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  dirty_1_15 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  dirty_1_16 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  dirty_1_17 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  dirty_1_18 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  dirty_1_19 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  dirty_1_20 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  dirty_1_21 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  dirty_1_22 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  dirty_1_23 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  dirty_1_24 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  dirty_1_25 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  dirty_1_26 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  dirty_1_27 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  dirty_1_28 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  dirty_1_29 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  dirty_1_30 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  dirty_1_31 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  dirty_1_32 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  dirty_1_33 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  dirty_1_34 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  dirty_1_35 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  dirty_1_36 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  dirty_1_37 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  dirty_1_38 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  dirty_1_39 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  dirty_1_40 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  dirty_1_41 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  dirty_1_42 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  dirty_1_43 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  dirty_1_44 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  dirty_1_45 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  dirty_1_46 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  dirty_1_47 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  dirty_1_48 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  dirty_1_49 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  dirty_1_50 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  dirty_1_51 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  dirty_1_52 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  dirty_1_53 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  dirty_1_54 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  dirty_1_55 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  dirty_1_56 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  dirty_1_57 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  dirty_1_58 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  dirty_1_59 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  dirty_1_60 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  dirty_1_61 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  dirty_1_62 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  dirty_1_63 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  dirty_1_64 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  dirty_1_65 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  dirty_1_66 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  dirty_1_67 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  dirty_1_68 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  dirty_1_69 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  dirty_1_70 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  dirty_1_71 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  dirty_1_72 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  dirty_1_73 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  dirty_1_74 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  dirty_1_75 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  dirty_1_76 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  dirty_1_77 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  dirty_1_78 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  dirty_1_79 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  dirty_1_80 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  dirty_1_81 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  dirty_1_82 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  dirty_1_83 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  dirty_1_84 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  dirty_1_85 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  dirty_1_86 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  dirty_1_87 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  dirty_1_88 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  dirty_1_89 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  dirty_1_90 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  dirty_1_91 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  dirty_1_92 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  dirty_1_93 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  dirty_1_94 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  dirty_1_95 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  dirty_1_96 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  dirty_1_97 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  dirty_1_98 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  dirty_1_99 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  dirty_1_100 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  dirty_1_101 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  dirty_1_102 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  dirty_1_103 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  dirty_1_104 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  dirty_1_105 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  dirty_1_106 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  dirty_1_107 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  dirty_1_108 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  dirty_1_109 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  dirty_1_110 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  dirty_1_111 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  dirty_1_112 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  dirty_1_113 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  dirty_1_114 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  dirty_1_115 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  dirty_1_116 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  dirty_1_117 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  dirty_1_118 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  dirty_1_119 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  dirty_1_120 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  dirty_1_121 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  dirty_1_122 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  dirty_1_123 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  dirty_1_124 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  dirty_1_125 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  dirty_1_126 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  dirty_1_127 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  dirty_1_128 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  dirty_1_129 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  dirty_1_130 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  dirty_1_131 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  dirty_1_132 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  dirty_1_133 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  dirty_1_134 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  dirty_1_135 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  dirty_1_136 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  dirty_1_137 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  dirty_1_138 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  dirty_1_139 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  dirty_1_140 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  dirty_1_141 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  dirty_1_142 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  dirty_1_143 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  dirty_1_144 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  dirty_1_145 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  dirty_1_146 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  dirty_1_147 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  dirty_1_148 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  dirty_1_149 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  dirty_1_150 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  dirty_1_151 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  dirty_1_152 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  dirty_1_153 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  dirty_1_154 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  dirty_1_155 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  dirty_1_156 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  dirty_1_157 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  dirty_1_158 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  dirty_1_159 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  dirty_1_160 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  dirty_1_161 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  dirty_1_162 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  dirty_1_163 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  dirty_1_164 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  dirty_1_165 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  dirty_1_166 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  dirty_1_167 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  dirty_1_168 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  dirty_1_169 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  dirty_1_170 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  dirty_1_171 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  dirty_1_172 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  dirty_1_173 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  dirty_1_174 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  dirty_1_175 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  dirty_1_176 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  dirty_1_177 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  dirty_1_178 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  dirty_1_179 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  dirty_1_180 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  dirty_1_181 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  dirty_1_182 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  dirty_1_183 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  dirty_1_184 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  dirty_1_185 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  dirty_1_186 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  dirty_1_187 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  dirty_1_188 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  dirty_1_189 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  dirty_1_190 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  dirty_1_191 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  dirty_1_192 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  dirty_1_193 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  dirty_1_194 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  dirty_1_195 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  dirty_1_196 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  dirty_1_197 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  dirty_1_198 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  dirty_1_199 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  dirty_1_200 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  dirty_1_201 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  dirty_1_202 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  dirty_1_203 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  dirty_1_204 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  dirty_1_205 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  dirty_1_206 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  dirty_1_207 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  dirty_1_208 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  dirty_1_209 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  dirty_1_210 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  dirty_1_211 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  dirty_1_212 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  dirty_1_213 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  dirty_1_214 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  dirty_1_215 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  dirty_1_216 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  dirty_1_217 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  dirty_1_218 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  dirty_1_219 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  dirty_1_220 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  dirty_1_221 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  dirty_1_222 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  dirty_1_223 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  dirty_1_224 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  dirty_1_225 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  dirty_1_226 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  dirty_1_227 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  dirty_1_228 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  dirty_1_229 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  dirty_1_230 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  dirty_1_231 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  dirty_1_232 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  dirty_1_233 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  dirty_1_234 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  dirty_1_235 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  dirty_1_236 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  dirty_1_237 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  dirty_1_238 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  dirty_1_239 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  dirty_1_240 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  dirty_1_241 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  dirty_1_242 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  dirty_1_243 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  dirty_1_244 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  dirty_1_245 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  dirty_1_246 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  dirty_1_247 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  dirty_1_248 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  dirty_1_249 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  dirty_1_250 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  dirty_1_251 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  dirty_1_252 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  dirty_1_253 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  dirty_1_254 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  dirty_1_255 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  req_valid = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  req_op = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  req_uncached = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  req_offset = _RAND_521[3:0];
  _RAND_522 = {1{`RANDOM}};
  req_lstype = _RAND_522[2:0];
  _RAND_523 = {1{`RANDOM}};
  req_set = _RAND_523[7:0];
  _RAND_524 = {1{`RANDOM}};
  req_tag = _RAND_524[19:0];
  _RAND_525 = {1{`RANDOM}};
  req_wstrb_0 = _RAND_525[3:0];
  _RAND_526 = {1{`RANDOM}};
  req_wdata_0 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  req_wdata_1 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  req_wstrb_1 = _RAND_528[3:0];
  _RAND_529 = {1{`RANDOM}};
  req_wline = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  req_wset = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  req_woffset = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  tagv_r_0 = _RAND_532[20:0];
  _RAND_533 = {1{`RANDOM}};
  tagv_r_1 = _RAND_533[20:0];
  _RAND_534 = {1{`RANDOM}};
  state = _RAND_534[2:0];
  _RAND_535 = {1{`RANDOM}};
  refillIDX_r = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  LFSR_result = _RAND_536[15:0];
  _RAND_537 = {1{`RANDOM}};
  wr_cnt = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  wstate = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  req_wline_1 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  req_woffset_1 = _RAND_540[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
